module SyncFifo(
  input        clock,
  input        reset,
  input        io_Writer_WriteEn, // @[src/main/scala/fifo_pkg/FifoPkg.scala 19:14]
  input  [8:0] io_Writer_WriteData, // @[src/main/scala/fifo_pkg/FifoPkg.scala 19:14]
  output       io_Writer_Full, // @[src/main/scala/fifo_pkg/FifoPkg.scala 19:14]
  input        io_Reader_ReadEn, // @[src/main/scala/fifo_pkg/FifoPkg.scala 19:14]
  output [8:0] io_Reader_ReadData, // @[src/main/scala/fifo_pkg/FifoPkg.scala 19:14]
  output       io_Reader_Empty // @[src/main/scala/fifo_pkg/FifoPkg.scala 19:14]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_198;
  reg [31:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [31:0] _RAND_201;
  reg [31:0] _RAND_202;
  reg [31:0] _RAND_203;
  reg [31:0] _RAND_204;
  reg [31:0] _RAND_205;
  reg [31:0] _RAND_206;
  reg [31:0] _RAND_207;
  reg [31:0] _RAND_208;
  reg [31:0] _RAND_209;
  reg [31:0] _RAND_210;
  reg [31:0] _RAND_211;
  reg [31:0] _RAND_212;
  reg [31:0] _RAND_213;
  reg [31:0] _RAND_214;
  reg [31:0] _RAND_215;
  reg [31:0] _RAND_216;
  reg [31:0] _RAND_217;
  reg [31:0] _RAND_218;
  reg [31:0] _RAND_219;
  reg [31:0] _RAND_220;
  reg [31:0] _RAND_221;
  reg [31:0] _RAND_222;
  reg [31:0] _RAND_223;
  reg [31:0] _RAND_224;
  reg [31:0] _RAND_225;
  reg [31:0] _RAND_226;
  reg [31:0] _RAND_227;
  reg [31:0] _RAND_228;
  reg [31:0] _RAND_229;
  reg [31:0] _RAND_230;
  reg [31:0] _RAND_231;
  reg [31:0] _RAND_232;
  reg [31:0] _RAND_233;
  reg [31:0] _RAND_234;
  reg [31:0] _RAND_235;
  reg [31:0] _RAND_236;
  reg [31:0] _RAND_237;
  reg [31:0] _RAND_238;
  reg [31:0] _RAND_239;
  reg [31:0] _RAND_240;
  reg [31:0] _RAND_241;
  reg [31:0] _RAND_242;
  reg [31:0] _RAND_243;
  reg [31:0] _RAND_244;
  reg [31:0] _RAND_245;
  reg [31:0] _RAND_246;
  reg [31:0] _RAND_247;
  reg [31:0] _RAND_248;
  reg [31:0] _RAND_249;
  reg [31:0] _RAND_250;
  reg [31:0] _RAND_251;
  reg [31:0] _RAND_252;
  reg [31:0] _RAND_253;
  reg [31:0] _RAND_254;
  reg [31:0] _RAND_255;
  reg [31:0] _RAND_256;
  reg [31:0] _RAND_257;
  reg [31:0] _RAND_258;
  reg [31:0] _RAND_259;
  reg [31:0] _RAND_260;
  reg [31:0] _RAND_261;
  reg [31:0] _RAND_262;
  reg [31:0] _RAND_263;
  reg [31:0] _RAND_264;
  reg [31:0] _RAND_265;
  reg [31:0] _RAND_266;
  reg [31:0] _RAND_267;
  reg [31:0] _RAND_268;
  reg [31:0] _RAND_269;
  reg [31:0] _RAND_270;
  reg [31:0] _RAND_271;
  reg [31:0] _RAND_272;
  reg [31:0] _RAND_273;
  reg [31:0] _RAND_274;
  reg [31:0] _RAND_275;
  reg [31:0] _RAND_276;
  reg [31:0] _RAND_277;
  reg [31:0] _RAND_278;
  reg [31:0] _RAND_279;
  reg [31:0] _RAND_280;
  reg [31:0] _RAND_281;
  reg [31:0] _RAND_282;
  reg [31:0] _RAND_283;
  reg [31:0] _RAND_284;
  reg [31:0] _RAND_285;
  reg [31:0] _RAND_286;
  reg [31:0] _RAND_287;
  reg [31:0] _RAND_288;
  reg [31:0] _RAND_289;
  reg [31:0] _RAND_290;
  reg [31:0] _RAND_291;
  reg [31:0] _RAND_292;
  reg [31:0] _RAND_293;
  reg [31:0] _RAND_294;
  reg [31:0] _RAND_295;
  reg [31:0] _RAND_296;
  reg [31:0] _RAND_297;
  reg [31:0] _RAND_298;
  reg [31:0] _RAND_299;
  reg [31:0] _RAND_300;
  reg [31:0] _RAND_301;
  reg [31:0] _RAND_302;
  reg [31:0] _RAND_303;
  reg [31:0] _RAND_304;
  reg [31:0] _RAND_305;
  reg [31:0] _RAND_306;
  reg [31:0] _RAND_307;
  reg [31:0] _RAND_308;
  reg [31:0] _RAND_309;
  reg [31:0] _RAND_310;
  reg [31:0] _RAND_311;
  reg [31:0] _RAND_312;
  reg [31:0] _RAND_313;
  reg [31:0] _RAND_314;
  reg [31:0] _RAND_315;
  reg [31:0] _RAND_316;
  reg [31:0] _RAND_317;
  reg [31:0] _RAND_318;
  reg [31:0] _RAND_319;
  reg [31:0] _RAND_320;
  reg [31:0] _RAND_321;
  reg [31:0] _RAND_322;
  reg [31:0] _RAND_323;
  reg [31:0] _RAND_324;
  reg [31:0] _RAND_325;
  reg [31:0] _RAND_326;
  reg [31:0] _RAND_327;
  reg [31:0] _RAND_328;
  reg [31:0] _RAND_329;
  reg [31:0] _RAND_330;
  reg [31:0] _RAND_331;
  reg [31:0] _RAND_332;
  reg [31:0] _RAND_333;
  reg [31:0] _RAND_334;
  reg [31:0] _RAND_335;
  reg [31:0] _RAND_336;
  reg [31:0] _RAND_337;
  reg [31:0] _RAND_338;
  reg [31:0] _RAND_339;
  reg [31:0] _RAND_340;
  reg [31:0] _RAND_341;
  reg [31:0] _RAND_342;
  reg [31:0] _RAND_343;
  reg [31:0] _RAND_344;
  reg [31:0] _RAND_345;
  reg [31:0] _RAND_346;
  reg [31:0] _RAND_347;
  reg [31:0] _RAND_348;
  reg [31:0] _RAND_349;
  reg [31:0] _RAND_350;
  reg [31:0] _RAND_351;
  reg [31:0] _RAND_352;
  reg [31:0] _RAND_353;
  reg [31:0] _RAND_354;
  reg [31:0] _RAND_355;
  reg [31:0] _RAND_356;
  reg [31:0] _RAND_357;
  reg [31:0] _RAND_358;
  reg [31:0] _RAND_359;
  reg [31:0] _RAND_360;
  reg [31:0] _RAND_361;
  reg [31:0] _RAND_362;
  reg [31:0] _RAND_363;
  reg [31:0] _RAND_364;
  reg [31:0] _RAND_365;
  reg [31:0] _RAND_366;
  reg [31:0] _RAND_367;
  reg [31:0] _RAND_368;
  reg [31:0] _RAND_369;
  reg [31:0] _RAND_370;
  reg [31:0] _RAND_371;
  reg [31:0] _RAND_372;
  reg [31:0] _RAND_373;
  reg [31:0] _RAND_374;
  reg [31:0] _RAND_375;
  reg [31:0] _RAND_376;
  reg [31:0] _RAND_377;
  reg [31:0] _RAND_378;
  reg [31:0] _RAND_379;
  reg [31:0] _RAND_380;
  reg [31:0] _RAND_381;
  reg [31:0] _RAND_382;
  reg [31:0] _RAND_383;
  reg [31:0] _RAND_384;
  reg [31:0] _RAND_385;
  reg [31:0] _RAND_386;
  reg [31:0] _RAND_387;
  reg [31:0] _RAND_388;
  reg [31:0] _RAND_389;
  reg [31:0] _RAND_390;
  reg [31:0] _RAND_391;
  reg [31:0] _RAND_392;
  reg [31:0] _RAND_393;
  reg [31:0] _RAND_394;
  reg [31:0] _RAND_395;
  reg [31:0] _RAND_396;
  reg [31:0] _RAND_397;
  reg [31:0] _RAND_398;
  reg [31:0] _RAND_399;
  reg [31:0] _RAND_400;
  reg [31:0] _RAND_401;
  reg [31:0] _RAND_402;
  reg [31:0] _RAND_403;
  reg [31:0] _RAND_404;
  reg [31:0] _RAND_405;
  reg [31:0] _RAND_406;
  reg [31:0] _RAND_407;
  reg [31:0] _RAND_408;
  reg [31:0] _RAND_409;
  reg [31:0] _RAND_410;
  reg [31:0] _RAND_411;
  reg [31:0] _RAND_412;
  reg [31:0] _RAND_413;
  reg [31:0] _RAND_414;
  reg [31:0] _RAND_415;
  reg [31:0] _RAND_416;
  reg [31:0] _RAND_417;
  reg [31:0] _RAND_418;
  reg [31:0] _RAND_419;
  reg [31:0] _RAND_420;
  reg [31:0] _RAND_421;
  reg [31:0] _RAND_422;
  reg [31:0] _RAND_423;
  reg [31:0] _RAND_424;
  reg [31:0] _RAND_425;
  reg [31:0] _RAND_426;
  reg [31:0] _RAND_427;
  reg [31:0] _RAND_428;
  reg [31:0] _RAND_429;
  reg [31:0] _RAND_430;
  reg [31:0] _RAND_431;
  reg [31:0] _RAND_432;
  reg [31:0] _RAND_433;
  reg [31:0] _RAND_434;
  reg [31:0] _RAND_435;
  reg [31:0] _RAND_436;
  reg [31:0] _RAND_437;
  reg [31:0] _RAND_438;
  reg [31:0] _RAND_439;
  reg [31:0] _RAND_440;
  reg [31:0] _RAND_441;
  reg [31:0] _RAND_442;
  reg [31:0] _RAND_443;
  reg [31:0] _RAND_444;
  reg [31:0] _RAND_445;
  reg [31:0] _RAND_446;
  reg [31:0] _RAND_447;
  reg [31:0] _RAND_448;
  reg [31:0] _RAND_449;
  reg [31:0] _RAND_450;
  reg [31:0] _RAND_451;
  reg [31:0] _RAND_452;
  reg [31:0] _RAND_453;
  reg [31:0] _RAND_454;
  reg [31:0] _RAND_455;
  reg [31:0] _RAND_456;
  reg [31:0] _RAND_457;
  reg [31:0] _RAND_458;
  reg [31:0] _RAND_459;
  reg [31:0] _RAND_460;
  reg [31:0] _RAND_461;
  reg [31:0] _RAND_462;
  reg [31:0] _RAND_463;
  reg [31:0] _RAND_464;
  reg [31:0] _RAND_465;
  reg [31:0] _RAND_466;
  reg [31:0] _RAND_467;
  reg [31:0] _RAND_468;
  reg [31:0] _RAND_469;
  reg [31:0] _RAND_470;
  reg [31:0] _RAND_471;
  reg [31:0] _RAND_472;
  reg [31:0] _RAND_473;
  reg [31:0] _RAND_474;
  reg [31:0] _RAND_475;
  reg [31:0] _RAND_476;
  reg [31:0] _RAND_477;
  reg [31:0] _RAND_478;
  reg [31:0] _RAND_479;
  reg [31:0] _RAND_480;
  reg [31:0] _RAND_481;
  reg [31:0] _RAND_482;
  reg [31:0] _RAND_483;
  reg [31:0] _RAND_484;
  reg [31:0] _RAND_485;
  reg [31:0] _RAND_486;
  reg [31:0] _RAND_487;
  reg [31:0] _RAND_488;
  reg [31:0] _RAND_489;
  reg [31:0] _RAND_490;
  reg [31:0] _RAND_491;
  reg [31:0] _RAND_492;
  reg [31:0] _RAND_493;
  reg [31:0] _RAND_494;
  reg [31:0] _RAND_495;
  reg [31:0] _RAND_496;
  reg [31:0] _RAND_497;
  reg [31:0] _RAND_498;
  reg [31:0] _RAND_499;
  reg [31:0] _RAND_500;
  reg [31:0] _RAND_501;
  reg [31:0] _RAND_502;
  reg [31:0] _RAND_503;
  reg [31:0] _RAND_504;
  reg [31:0] _RAND_505;
  reg [31:0] _RAND_506;
  reg [31:0] _RAND_507;
  reg [31:0] _RAND_508;
  reg [31:0] _RAND_509;
  reg [31:0] _RAND_510;
  reg [31:0] _RAND_511;
  reg [31:0] _RAND_512;
  reg [31:0] _RAND_513;
  reg [31:0] _RAND_514;
  reg [31:0] _RAND_515;
  reg [31:0] _RAND_516;
  reg [31:0] _RAND_517;
  reg [31:0] _RAND_518;
  reg [31:0] _RAND_519;
  reg [31:0] _RAND_520;
  reg [31:0] _RAND_521;
  reg [31:0] _RAND_522;
  reg [31:0] _RAND_523;
  reg [31:0] _RAND_524;
  reg [31:0] _RAND_525;
  reg [31:0] _RAND_526;
  reg [31:0] _RAND_527;
  reg [31:0] _RAND_528;
  reg [31:0] _RAND_529;
  reg [31:0] _RAND_530;
  reg [31:0] _RAND_531;
  reg [31:0] _RAND_532;
  reg [31:0] _RAND_533;
  reg [31:0] _RAND_534;
  reg [31:0] _RAND_535;
  reg [31:0] _RAND_536;
  reg [31:0] _RAND_537;
  reg [31:0] _RAND_538;
  reg [31:0] _RAND_539;
  reg [31:0] _RAND_540;
  reg [31:0] _RAND_541;
  reg [31:0] _RAND_542;
  reg [31:0] _RAND_543;
  reg [31:0] _RAND_544;
  reg [31:0] _RAND_545;
  reg [31:0] _RAND_546;
  reg [31:0] _RAND_547;
  reg [31:0] _RAND_548;
  reg [31:0] _RAND_549;
  reg [31:0] _RAND_550;
  reg [31:0] _RAND_551;
  reg [31:0] _RAND_552;
  reg [31:0] _RAND_553;
  reg [31:0] _RAND_554;
  reg [31:0] _RAND_555;
  reg [31:0] _RAND_556;
  reg [31:0] _RAND_557;
  reg [31:0] _RAND_558;
  reg [31:0] _RAND_559;
  reg [31:0] _RAND_560;
  reg [31:0] _RAND_561;
  reg [31:0] _RAND_562;
  reg [31:0] _RAND_563;
  reg [31:0] _RAND_564;
  reg [31:0] _RAND_565;
  reg [31:0] _RAND_566;
  reg [31:0] _RAND_567;
  reg [31:0] _RAND_568;
  reg [31:0] _RAND_569;
  reg [31:0] _RAND_570;
  reg [31:0] _RAND_571;
  reg [31:0] _RAND_572;
  reg [31:0] _RAND_573;
  reg [31:0] _RAND_574;
  reg [31:0] _RAND_575;
  reg [31:0] _RAND_576;
  reg [31:0] _RAND_577;
  reg [31:0] _RAND_578;
  reg [31:0] _RAND_579;
  reg [31:0] _RAND_580;
  reg [31:0] _RAND_581;
  reg [31:0] _RAND_582;
  reg [31:0] _RAND_583;
  reg [31:0] _RAND_584;
  reg [31:0] _RAND_585;
  reg [31:0] _RAND_586;
  reg [31:0] _RAND_587;
  reg [31:0] _RAND_588;
  reg [31:0] _RAND_589;
  reg [31:0] _RAND_590;
  reg [31:0] _RAND_591;
  reg [31:0] _RAND_592;
  reg [31:0] _RAND_593;
  reg [31:0] _RAND_594;
  reg [31:0] _RAND_595;
  reg [31:0] _RAND_596;
  reg [31:0] _RAND_597;
  reg [31:0] _RAND_598;
  reg [31:0] _RAND_599;
  reg [31:0] _RAND_600;
  reg [31:0] _RAND_601;
  reg [31:0] _RAND_602;
  reg [31:0] _RAND_603;
  reg [31:0] _RAND_604;
  reg [31:0] _RAND_605;
  reg [31:0] _RAND_606;
  reg [31:0] _RAND_607;
  reg [31:0] _RAND_608;
  reg [31:0] _RAND_609;
  reg [31:0] _RAND_610;
  reg [31:0] _RAND_611;
  reg [31:0] _RAND_612;
  reg [31:0] _RAND_613;
  reg [31:0] _RAND_614;
  reg [31:0] _RAND_615;
  reg [31:0] _RAND_616;
  reg [31:0] _RAND_617;
  reg [31:0] _RAND_618;
  reg [31:0] _RAND_619;
  reg [31:0] _RAND_620;
  reg [31:0] _RAND_621;
  reg [31:0] _RAND_622;
  reg [31:0] _RAND_623;
  reg [31:0] _RAND_624;
  reg [31:0] _RAND_625;
  reg [31:0] _RAND_626;
  reg [31:0] _RAND_627;
  reg [31:0] _RAND_628;
  reg [31:0] _RAND_629;
  reg [31:0] _RAND_630;
  reg [31:0] _RAND_631;
  reg [31:0] _RAND_632;
  reg [31:0] _RAND_633;
  reg [31:0] _RAND_634;
  reg [31:0] _RAND_635;
  reg [31:0] _RAND_636;
  reg [31:0] _RAND_637;
  reg [31:0] _RAND_638;
  reg [31:0] _RAND_639;
  reg [31:0] _RAND_640;
  reg [31:0] _RAND_641;
  reg [31:0] _RAND_642;
  reg [31:0] _RAND_643;
  reg [31:0] _RAND_644;
  reg [31:0] _RAND_645;
  reg [31:0] _RAND_646;
  reg [31:0] _RAND_647;
  reg [31:0] _RAND_648;
  reg [31:0] _RAND_649;
  reg [31:0] _RAND_650;
  reg [31:0] _RAND_651;
  reg [31:0] _RAND_652;
  reg [31:0] _RAND_653;
  reg [31:0] _RAND_654;
  reg [31:0] _RAND_655;
  reg [31:0] _RAND_656;
  reg [31:0] _RAND_657;
  reg [31:0] _RAND_658;
  reg [31:0] _RAND_659;
  reg [31:0] _RAND_660;
  reg [31:0] _RAND_661;
  reg [31:0] _RAND_662;
  reg [31:0] _RAND_663;
  reg [31:0] _RAND_664;
  reg [31:0] _RAND_665;
  reg [31:0] _RAND_666;
  reg [31:0] _RAND_667;
  reg [31:0] _RAND_668;
  reg [31:0] _RAND_669;
  reg [31:0] _RAND_670;
  reg [31:0] _RAND_671;
  reg [31:0] _RAND_672;
  reg [31:0] _RAND_673;
  reg [31:0] _RAND_674;
  reg [31:0] _RAND_675;
  reg [31:0] _RAND_676;
  reg [31:0] _RAND_677;
  reg [31:0] _RAND_678;
  reg [31:0] _RAND_679;
  reg [31:0] _RAND_680;
  reg [31:0] _RAND_681;
  reg [31:0] _RAND_682;
  reg [31:0] _RAND_683;
  reg [31:0] _RAND_684;
  reg [31:0] _RAND_685;
  reg [31:0] _RAND_686;
  reg [31:0] _RAND_687;
  reg [31:0] _RAND_688;
  reg [31:0] _RAND_689;
  reg [31:0] _RAND_690;
  reg [31:0] _RAND_691;
  reg [31:0] _RAND_692;
  reg [31:0] _RAND_693;
  reg [31:0] _RAND_694;
  reg [31:0] _RAND_695;
  reg [31:0] _RAND_696;
  reg [31:0] _RAND_697;
  reg [31:0] _RAND_698;
  reg [31:0] _RAND_699;
  reg [31:0] _RAND_700;
  reg [31:0] _RAND_701;
  reg [31:0] _RAND_702;
  reg [31:0] _RAND_703;
  reg [31:0] _RAND_704;
  reg [31:0] _RAND_705;
  reg [31:0] _RAND_706;
  reg [31:0] _RAND_707;
  reg [31:0] _RAND_708;
  reg [31:0] _RAND_709;
  reg [31:0] _RAND_710;
  reg [31:0] _RAND_711;
  reg [31:0] _RAND_712;
  reg [31:0] _RAND_713;
  reg [31:0] _RAND_714;
  reg [31:0] _RAND_715;
  reg [31:0] _RAND_716;
  reg [31:0] _RAND_717;
  reg [31:0] _RAND_718;
  reg [31:0] _RAND_719;
  reg [31:0] _RAND_720;
  reg [31:0] _RAND_721;
  reg [31:0] _RAND_722;
  reg [31:0] _RAND_723;
  reg [31:0] _RAND_724;
  reg [31:0] _RAND_725;
  reg [31:0] _RAND_726;
  reg [31:0] _RAND_727;
  reg [31:0] _RAND_728;
  reg [31:0] _RAND_729;
  reg [31:0] _RAND_730;
  reg [31:0] _RAND_731;
  reg [31:0] _RAND_732;
  reg [31:0] _RAND_733;
  reg [31:0] _RAND_734;
  reg [31:0] _RAND_735;
  reg [31:0] _RAND_736;
  reg [31:0] _RAND_737;
  reg [31:0] _RAND_738;
  reg [31:0] _RAND_739;
  reg [31:0] _RAND_740;
  reg [31:0] _RAND_741;
  reg [31:0] _RAND_742;
  reg [31:0] _RAND_743;
  reg [31:0] _RAND_744;
  reg [31:0] _RAND_745;
  reg [31:0] _RAND_746;
  reg [31:0] _RAND_747;
  reg [31:0] _RAND_748;
  reg [31:0] _RAND_749;
  reg [31:0] _RAND_750;
  reg [31:0] _RAND_751;
  reg [31:0] _RAND_752;
  reg [31:0] _RAND_753;
  reg [31:0] _RAND_754;
  reg [31:0] _RAND_755;
  reg [31:0] _RAND_756;
  reg [31:0] _RAND_757;
  reg [31:0] _RAND_758;
  reg [31:0] _RAND_759;
  reg [31:0] _RAND_760;
  reg [31:0] _RAND_761;
  reg [31:0] _RAND_762;
  reg [31:0] _RAND_763;
  reg [31:0] _RAND_764;
  reg [31:0] _RAND_765;
  reg [31:0] _RAND_766;
  reg [31:0] _RAND_767;
  reg [31:0] _RAND_768;
  reg [31:0] _RAND_769;
  reg [31:0] _RAND_770;
  reg [31:0] _RAND_771;
  reg [31:0] _RAND_772;
  reg [31:0] _RAND_773;
  reg [31:0] _RAND_774;
  reg [31:0] _RAND_775;
  reg [31:0] _RAND_776;
  reg [31:0] _RAND_777;
  reg [31:0] _RAND_778;
  reg [31:0] _RAND_779;
  reg [31:0] _RAND_780;
  reg [31:0] _RAND_781;
  reg [31:0] _RAND_782;
  reg [31:0] _RAND_783;
  reg [31:0] _RAND_784;
  reg [31:0] _RAND_785;
  reg [31:0] _RAND_786;
  reg [31:0] _RAND_787;
  reg [31:0] _RAND_788;
  reg [31:0] _RAND_789;
  reg [31:0] _RAND_790;
  reg [31:0] _RAND_791;
  reg [31:0] _RAND_792;
  reg [31:0] _RAND_793;
  reg [31:0] _RAND_794;
  reg [31:0] _RAND_795;
  reg [31:0] _RAND_796;
  reg [31:0] _RAND_797;
  reg [31:0] _RAND_798;
  reg [31:0] _RAND_799;
  reg [31:0] _RAND_800;
  reg [31:0] _RAND_801;
  reg [31:0] _RAND_802;
  reg [31:0] _RAND_803;
  reg [31:0] _RAND_804;
  reg [31:0] _RAND_805;
  reg [31:0] _RAND_806;
  reg [31:0] _RAND_807;
  reg [31:0] _RAND_808;
  reg [31:0] _RAND_809;
  reg [31:0] _RAND_810;
  reg [31:0] _RAND_811;
  reg [31:0] _RAND_812;
  reg [31:0] _RAND_813;
  reg [31:0] _RAND_814;
  reg [31:0] _RAND_815;
  reg [31:0] _RAND_816;
  reg [31:0] _RAND_817;
  reg [31:0] _RAND_818;
  reg [31:0] _RAND_819;
  reg [31:0] _RAND_820;
  reg [31:0] _RAND_821;
  reg [31:0] _RAND_822;
  reg [31:0] _RAND_823;
  reg [31:0] _RAND_824;
  reg [31:0] _RAND_825;
  reg [31:0] _RAND_826;
  reg [31:0] _RAND_827;
  reg [31:0] _RAND_828;
  reg [31:0] _RAND_829;
  reg [31:0] _RAND_830;
  reg [31:0] _RAND_831;
  reg [31:0] _RAND_832;
  reg [31:0] _RAND_833;
  reg [31:0] _RAND_834;
  reg [31:0] _RAND_835;
  reg [31:0] _RAND_836;
  reg [31:0] _RAND_837;
  reg [31:0] _RAND_838;
  reg [31:0] _RAND_839;
  reg [31:0] _RAND_840;
  reg [31:0] _RAND_841;
  reg [31:0] _RAND_842;
  reg [31:0] _RAND_843;
  reg [31:0] _RAND_844;
  reg [31:0] _RAND_845;
  reg [31:0] _RAND_846;
  reg [31:0] _RAND_847;
  reg [31:0] _RAND_848;
  reg [31:0] _RAND_849;
  reg [31:0] _RAND_850;
  reg [31:0] _RAND_851;
  reg [31:0] _RAND_852;
  reg [31:0] _RAND_853;
  reg [31:0] _RAND_854;
  reg [31:0] _RAND_855;
  reg [31:0] _RAND_856;
  reg [31:0] _RAND_857;
  reg [31:0] _RAND_858;
  reg [31:0] _RAND_859;
  reg [31:0] _RAND_860;
  reg [31:0] _RAND_861;
  reg [31:0] _RAND_862;
  reg [31:0] _RAND_863;
  reg [31:0] _RAND_864;
  reg [31:0] _RAND_865;
  reg [31:0] _RAND_866;
  reg [31:0] _RAND_867;
  reg [31:0] _RAND_868;
  reg [31:0] _RAND_869;
  reg [31:0] _RAND_870;
  reg [31:0] _RAND_871;
  reg [31:0] _RAND_872;
  reg [31:0] _RAND_873;
  reg [31:0] _RAND_874;
  reg [31:0] _RAND_875;
  reg [31:0] _RAND_876;
  reg [31:0] _RAND_877;
  reg [31:0] _RAND_878;
  reg [31:0] _RAND_879;
  reg [31:0] _RAND_880;
  reg [31:0] _RAND_881;
  reg [31:0] _RAND_882;
  reg [31:0] _RAND_883;
  reg [31:0] _RAND_884;
  reg [31:0] _RAND_885;
  reg [31:0] _RAND_886;
  reg [31:0] _RAND_887;
  reg [31:0] _RAND_888;
  reg [31:0] _RAND_889;
  reg [31:0] _RAND_890;
  reg [31:0] _RAND_891;
  reg [31:0] _RAND_892;
  reg [31:0] _RAND_893;
  reg [31:0] _RAND_894;
  reg [31:0] _RAND_895;
  reg [31:0] _RAND_896;
  reg [31:0] _RAND_897;
  reg [31:0] _RAND_898;
  reg [31:0] _RAND_899;
  reg [31:0] _RAND_900;
  reg [31:0] _RAND_901;
  reg [31:0] _RAND_902;
  reg [31:0] _RAND_903;
  reg [31:0] _RAND_904;
  reg [31:0] _RAND_905;
  reg [31:0] _RAND_906;
  reg [31:0] _RAND_907;
  reg [31:0] _RAND_908;
  reg [31:0] _RAND_909;
  reg [31:0] _RAND_910;
  reg [31:0] _RAND_911;
  reg [31:0] _RAND_912;
  reg [31:0] _RAND_913;
  reg [31:0] _RAND_914;
  reg [31:0] _RAND_915;
  reg [31:0] _RAND_916;
  reg [31:0] _RAND_917;
  reg [31:0] _RAND_918;
  reg [31:0] _RAND_919;
  reg [31:0] _RAND_920;
  reg [31:0] _RAND_921;
  reg [31:0] _RAND_922;
  reg [31:0] _RAND_923;
  reg [31:0] _RAND_924;
  reg [31:0] _RAND_925;
  reg [31:0] _RAND_926;
  reg [31:0] _RAND_927;
  reg [31:0] _RAND_928;
  reg [31:0] _RAND_929;
  reg [31:0] _RAND_930;
  reg [31:0] _RAND_931;
  reg [31:0] _RAND_932;
  reg [31:0] _RAND_933;
  reg [31:0] _RAND_934;
  reg [31:0] _RAND_935;
  reg [31:0] _RAND_936;
  reg [31:0] _RAND_937;
  reg [31:0] _RAND_938;
  reg [31:0] _RAND_939;
  reg [31:0] _RAND_940;
  reg [31:0] _RAND_941;
  reg [31:0] _RAND_942;
  reg [31:0] _RAND_943;
  reg [31:0] _RAND_944;
  reg [31:0] _RAND_945;
  reg [31:0] _RAND_946;
  reg [31:0] _RAND_947;
  reg [31:0] _RAND_948;
  reg [31:0] _RAND_949;
  reg [31:0] _RAND_950;
  reg [31:0] _RAND_951;
  reg [31:0] _RAND_952;
  reg [31:0] _RAND_953;
  reg [31:0] _RAND_954;
  reg [31:0] _RAND_955;
  reg [31:0] _RAND_956;
  reg [31:0] _RAND_957;
  reg [31:0] _RAND_958;
  reg [31:0] _RAND_959;
  reg [31:0] _RAND_960;
  reg [31:0] _RAND_961;
  reg [31:0] _RAND_962;
  reg [31:0] _RAND_963;
  reg [31:0] _RAND_964;
  reg [31:0] _RAND_965;
  reg [31:0] _RAND_966;
  reg [31:0] _RAND_967;
  reg [31:0] _RAND_968;
  reg [31:0] _RAND_969;
  reg [31:0] _RAND_970;
  reg [31:0] _RAND_971;
  reg [31:0] _RAND_972;
  reg [31:0] _RAND_973;
  reg [31:0] _RAND_974;
  reg [31:0] _RAND_975;
  reg [31:0] _RAND_976;
  reg [31:0] _RAND_977;
  reg [31:0] _RAND_978;
  reg [31:0] _RAND_979;
  reg [31:0] _RAND_980;
  reg [31:0] _RAND_981;
  reg [31:0] _RAND_982;
  reg [31:0] _RAND_983;
  reg [31:0] _RAND_984;
  reg [31:0] _RAND_985;
  reg [31:0] _RAND_986;
  reg [31:0] _RAND_987;
  reg [31:0] _RAND_988;
  reg [31:0] _RAND_989;
  reg [31:0] _RAND_990;
  reg [31:0] _RAND_991;
  reg [31:0] _RAND_992;
  reg [31:0] _RAND_993;
  reg [31:0] _RAND_994;
  reg [31:0] _RAND_995;
  reg [31:0] _RAND_996;
  reg [31:0] _RAND_997;
  reg [31:0] _RAND_998;
  reg [31:0] _RAND_999;
  reg [31:0] _RAND_1000;
  reg [31:0] _RAND_1001;
  reg [31:0] _RAND_1002;
  reg [31:0] _RAND_1003;
  reg [31:0] _RAND_1004;
  reg [31:0] _RAND_1005;
  reg [31:0] _RAND_1006;
  reg [31:0] _RAND_1007;
  reg [31:0] _RAND_1008;
  reg [31:0] _RAND_1009;
  reg [31:0] _RAND_1010;
  reg [31:0] _RAND_1011;
  reg [31:0] _RAND_1012;
  reg [31:0] _RAND_1013;
  reg [31:0] _RAND_1014;
  reg [31:0] _RAND_1015;
  reg [31:0] _RAND_1016;
  reg [31:0] _RAND_1017;
  reg [31:0] _RAND_1018;
  reg [31:0] _RAND_1019;
  reg [31:0] _RAND_1020;
  reg [31:0] _RAND_1021;
  reg [31:0] _RAND_1022;
  reg [31:0] _RAND_1023;
  reg [31:0] _RAND_1024;
  reg [31:0] _RAND_1025;
`endif // RANDOMIZE_REG_INIT
  reg [10:0] WritePtr; // @[src/main/scala/fifo_pkg/FifoPkg.scala 26:25]
  reg [10:0] ReadPtr; // @[src/main/scala/fifo_pkg/FifoPkg.scala 27:24]
  reg [8:0] FifoCell_0; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_1; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_2; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_3; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_4; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_5; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_6; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_7; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_8; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_9; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_10; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_11; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_12; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_13; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_14; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_15; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_16; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_17; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_18; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_19; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_20; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_21; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_22; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_23; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_24; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_25; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_26; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_27; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_28; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_29; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_30; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_31; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_32; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_33; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_34; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_35; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_36; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_37; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_38; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_39; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_40; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_41; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_42; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_43; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_44; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_45; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_46; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_47; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_48; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_49; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_50; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_51; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_52; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_53; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_54; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_55; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_56; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_57; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_58; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_59; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_60; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_61; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_62; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_63; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_64; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_65; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_66; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_67; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_68; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_69; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_70; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_71; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_72; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_73; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_74; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_75; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_76; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_77; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_78; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_79; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_80; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_81; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_82; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_83; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_84; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_85; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_86; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_87; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_88; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_89; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_90; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_91; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_92; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_93; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_94; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_95; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_96; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_97; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_98; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_99; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_100; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_101; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_102; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_103; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_104; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_105; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_106; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_107; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_108; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_109; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_110; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_111; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_112; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_113; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_114; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_115; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_116; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_117; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_118; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_119; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_120; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_121; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_122; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_123; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_124; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_125; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_126; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_127; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_128; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_129; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_130; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_131; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_132; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_133; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_134; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_135; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_136; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_137; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_138; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_139; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_140; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_141; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_142; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_143; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_144; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_145; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_146; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_147; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_148; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_149; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_150; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_151; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_152; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_153; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_154; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_155; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_156; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_157; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_158; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_159; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_160; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_161; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_162; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_163; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_164; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_165; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_166; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_167; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_168; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_169; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_170; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_171; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_172; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_173; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_174; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_175; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_176; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_177; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_178; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_179; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_180; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_181; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_182; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_183; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_184; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_185; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_186; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_187; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_188; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_189; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_190; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_191; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_192; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_193; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_194; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_195; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_196; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_197; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_198; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_199; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_200; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_201; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_202; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_203; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_204; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_205; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_206; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_207; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_208; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_209; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_210; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_211; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_212; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_213; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_214; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_215; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_216; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_217; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_218; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_219; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_220; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_221; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_222; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_223; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_224; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_225; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_226; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_227; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_228; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_229; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_230; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_231; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_232; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_233; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_234; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_235; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_236; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_237; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_238; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_239; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_240; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_241; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_242; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_243; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_244; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_245; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_246; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_247; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_248; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_249; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_250; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_251; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_252; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_253; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_254; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_255; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_256; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_257; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_258; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_259; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_260; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_261; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_262; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_263; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_264; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_265; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_266; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_267; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_268; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_269; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_270; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_271; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_272; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_273; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_274; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_275; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_276; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_277; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_278; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_279; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_280; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_281; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_282; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_283; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_284; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_285; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_286; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_287; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_288; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_289; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_290; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_291; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_292; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_293; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_294; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_295; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_296; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_297; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_298; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_299; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_300; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_301; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_302; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_303; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_304; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_305; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_306; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_307; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_308; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_309; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_310; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_311; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_312; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_313; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_314; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_315; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_316; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_317; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_318; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_319; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_320; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_321; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_322; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_323; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_324; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_325; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_326; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_327; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_328; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_329; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_330; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_331; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_332; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_333; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_334; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_335; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_336; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_337; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_338; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_339; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_340; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_341; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_342; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_343; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_344; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_345; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_346; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_347; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_348; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_349; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_350; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_351; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_352; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_353; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_354; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_355; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_356; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_357; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_358; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_359; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_360; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_361; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_362; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_363; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_364; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_365; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_366; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_367; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_368; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_369; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_370; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_371; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_372; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_373; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_374; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_375; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_376; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_377; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_378; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_379; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_380; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_381; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_382; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_383; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_384; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_385; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_386; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_387; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_388; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_389; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_390; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_391; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_392; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_393; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_394; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_395; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_396; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_397; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_398; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_399; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_400; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_401; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_402; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_403; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_404; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_405; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_406; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_407; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_408; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_409; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_410; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_411; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_412; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_413; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_414; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_415; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_416; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_417; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_418; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_419; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_420; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_421; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_422; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_423; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_424; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_425; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_426; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_427; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_428; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_429; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_430; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_431; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_432; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_433; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_434; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_435; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_436; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_437; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_438; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_439; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_440; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_441; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_442; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_443; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_444; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_445; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_446; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_447; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_448; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_449; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_450; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_451; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_452; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_453; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_454; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_455; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_456; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_457; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_458; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_459; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_460; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_461; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_462; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_463; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_464; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_465; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_466; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_467; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_468; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_469; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_470; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_471; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_472; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_473; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_474; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_475; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_476; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_477; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_478; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_479; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_480; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_481; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_482; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_483; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_484; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_485; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_486; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_487; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_488; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_489; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_490; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_491; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_492; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_493; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_494; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_495; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_496; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_497; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_498; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_499; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_500; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_501; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_502; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_503; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_504; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_505; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_506; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_507; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_508; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_509; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_510; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_511; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_512; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_513; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_514; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_515; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_516; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_517; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_518; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_519; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_520; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_521; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_522; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_523; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_524; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_525; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_526; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_527; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_528; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_529; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_530; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_531; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_532; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_533; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_534; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_535; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_536; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_537; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_538; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_539; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_540; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_541; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_542; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_543; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_544; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_545; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_546; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_547; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_548; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_549; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_550; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_551; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_552; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_553; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_554; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_555; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_556; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_557; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_558; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_559; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_560; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_561; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_562; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_563; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_564; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_565; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_566; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_567; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_568; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_569; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_570; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_571; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_572; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_573; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_574; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_575; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_576; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_577; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_578; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_579; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_580; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_581; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_582; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_583; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_584; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_585; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_586; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_587; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_588; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_589; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_590; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_591; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_592; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_593; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_594; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_595; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_596; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_597; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_598; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_599; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_600; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_601; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_602; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_603; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_604; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_605; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_606; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_607; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_608; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_609; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_610; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_611; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_612; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_613; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_614; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_615; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_616; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_617; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_618; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_619; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_620; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_621; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_622; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_623; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_624; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_625; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_626; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_627; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_628; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_629; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_630; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_631; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_632; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_633; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_634; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_635; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_636; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_637; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_638; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_639; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_640; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_641; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_642; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_643; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_644; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_645; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_646; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_647; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_648; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_649; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_650; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_651; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_652; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_653; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_654; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_655; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_656; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_657; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_658; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_659; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_660; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_661; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_662; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_663; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_664; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_665; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_666; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_667; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_668; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_669; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_670; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_671; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_672; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_673; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_674; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_675; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_676; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_677; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_678; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_679; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_680; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_681; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_682; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_683; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_684; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_685; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_686; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_687; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_688; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_689; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_690; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_691; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_692; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_693; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_694; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_695; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_696; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_697; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_698; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_699; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_700; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_701; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_702; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_703; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_704; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_705; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_706; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_707; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_708; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_709; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_710; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_711; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_712; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_713; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_714; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_715; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_716; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_717; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_718; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_719; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_720; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_721; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_722; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_723; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_724; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_725; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_726; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_727; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_728; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_729; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_730; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_731; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_732; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_733; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_734; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_735; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_736; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_737; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_738; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_739; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_740; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_741; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_742; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_743; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_744; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_745; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_746; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_747; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_748; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_749; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_750; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_751; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_752; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_753; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_754; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_755; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_756; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_757; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_758; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_759; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_760; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_761; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_762; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_763; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_764; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_765; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_766; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_767; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_768; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_769; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_770; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_771; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_772; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_773; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_774; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_775; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_776; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_777; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_778; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_779; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_780; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_781; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_782; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_783; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_784; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_785; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_786; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_787; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_788; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_789; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_790; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_791; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_792; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_793; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_794; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_795; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_796; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_797; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_798; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_799; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_800; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_801; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_802; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_803; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_804; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_805; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_806; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_807; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_808; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_809; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_810; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_811; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_812; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_813; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_814; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_815; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_816; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_817; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_818; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_819; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_820; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_821; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_822; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_823; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_824; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_825; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_826; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_827; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_828; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_829; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_830; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_831; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_832; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_833; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_834; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_835; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_836; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_837; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_838; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_839; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_840; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_841; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_842; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_843; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_844; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_845; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_846; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_847; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_848; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_849; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_850; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_851; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_852; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_853; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_854; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_855; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_856; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_857; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_858; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_859; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_860; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_861; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_862; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_863; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_864; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_865; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_866; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_867; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_868; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_869; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_870; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_871; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_872; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_873; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_874; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_875; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_876; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_877; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_878; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_879; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_880; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_881; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_882; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_883; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_884; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_885; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_886; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_887; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_888; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_889; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_890; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_891; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_892; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_893; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_894; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_895; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_896; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_897; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_898; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_899; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_900; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_901; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_902; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_903; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_904; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_905; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_906; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_907; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_908; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_909; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_910; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_911; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_912; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_913; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_914; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_915; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_916; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_917; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_918; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_919; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_920; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_921; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_922; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_923; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_924; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_925; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_926; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_927; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_928; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_929; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_930; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_931; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_932; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_933; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_934; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_935; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_936; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_937; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_938; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_939; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_940; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_941; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_942; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_943; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_944; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_945; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_946; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_947; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_948; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_949; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_950; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_951; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_952; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_953; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_954; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_955; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_956; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_957; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_958; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_959; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_960; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_961; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_962; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_963; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_964; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_965; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_966; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_967; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_968; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_969; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_970; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_971; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_972; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_973; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_974; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_975; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_976; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_977; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_978; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_979; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_980; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_981; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_982; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_983; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_984; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_985; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_986; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_987; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_988; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_989; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_990; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_991; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_992; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_993; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_994; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_995; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_996; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_997; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_998; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_999; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_1000; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_1001; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_1002; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_1003; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_1004; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_1005; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_1006; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_1007; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_1008; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_1009; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_1010; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_1011; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_1012; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_1013; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_1014; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_1015; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_1016; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_1017; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_1018; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_1019; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_1020; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_1021; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_1022; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  reg [8:0] FifoCell_1023; // @[src/main/scala/fifo_pkg/FifoPkg.scala 28:21]
  wire  _io_Writer_Full_T_5 = WritePtr[9:0] == ReadPtr[9:0]; // @[src/main/scala/fifo_pkg/FifoPkg.scala 31:54]
  wire  _T_2 = ~io_Writer_Full & io_Writer_WriteEn; // @[src/main/scala/fifo_pkg/FifoPkg.scala 34:32]
  wire [10:0] _WritePtr_T_1 = WritePtr + 11'h1; // @[src/main/scala/fifo_pkg/FifoPkg.scala 35:26]
  wire [10:0] _ReadPtr_T_1 = ReadPtr + 11'h1; // @[src/main/scala/fifo_pkg/FifoPkg.scala 39:24]
  wire [8:0] _GEN_2051 = 10'h1 == ReadPtr[9:0] ? FifoCell_1 : FifoCell_0; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2052 = 10'h2 == ReadPtr[9:0] ? FifoCell_2 : _GEN_2051; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2053 = 10'h3 == ReadPtr[9:0] ? FifoCell_3 : _GEN_2052; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2054 = 10'h4 == ReadPtr[9:0] ? FifoCell_4 : _GEN_2053; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2055 = 10'h5 == ReadPtr[9:0] ? FifoCell_5 : _GEN_2054; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2056 = 10'h6 == ReadPtr[9:0] ? FifoCell_6 : _GEN_2055; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2057 = 10'h7 == ReadPtr[9:0] ? FifoCell_7 : _GEN_2056; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2058 = 10'h8 == ReadPtr[9:0] ? FifoCell_8 : _GEN_2057; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2059 = 10'h9 == ReadPtr[9:0] ? FifoCell_9 : _GEN_2058; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2060 = 10'ha == ReadPtr[9:0] ? FifoCell_10 : _GEN_2059; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2061 = 10'hb == ReadPtr[9:0] ? FifoCell_11 : _GEN_2060; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2062 = 10'hc == ReadPtr[9:0] ? FifoCell_12 : _GEN_2061; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2063 = 10'hd == ReadPtr[9:0] ? FifoCell_13 : _GEN_2062; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2064 = 10'he == ReadPtr[9:0] ? FifoCell_14 : _GEN_2063; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2065 = 10'hf == ReadPtr[9:0] ? FifoCell_15 : _GEN_2064; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2066 = 10'h10 == ReadPtr[9:0] ? FifoCell_16 : _GEN_2065; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2067 = 10'h11 == ReadPtr[9:0] ? FifoCell_17 : _GEN_2066; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2068 = 10'h12 == ReadPtr[9:0] ? FifoCell_18 : _GEN_2067; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2069 = 10'h13 == ReadPtr[9:0] ? FifoCell_19 : _GEN_2068; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2070 = 10'h14 == ReadPtr[9:0] ? FifoCell_20 : _GEN_2069; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2071 = 10'h15 == ReadPtr[9:0] ? FifoCell_21 : _GEN_2070; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2072 = 10'h16 == ReadPtr[9:0] ? FifoCell_22 : _GEN_2071; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2073 = 10'h17 == ReadPtr[9:0] ? FifoCell_23 : _GEN_2072; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2074 = 10'h18 == ReadPtr[9:0] ? FifoCell_24 : _GEN_2073; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2075 = 10'h19 == ReadPtr[9:0] ? FifoCell_25 : _GEN_2074; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2076 = 10'h1a == ReadPtr[9:0] ? FifoCell_26 : _GEN_2075; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2077 = 10'h1b == ReadPtr[9:0] ? FifoCell_27 : _GEN_2076; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2078 = 10'h1c == ReadPtr[9:0] ? FifoCell_28 : _GEN_2077; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2079 = 10'h1d == ReadPtr[9:0] ? FifoCell_29 : _GEN_2078; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2080 = 10'h1e == ReadPtr[9:0] ? FifoCell_30 : _GEN_2079; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2081 = 10'h1f == ReadPtr[9:0] ? FifoCell_31 : _GEN_2080; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2082 = 10'h20 == ReadPtr[9:0] ? FifoCell_32 : _GEN_2081; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2083 = 10'h21 == ReadPtr[9:0] ? FifoCell_33 : _GEN_2082; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2084 = 10'h22 == ReadPtr[9:0] ? FifoCell_34 : _GEN_2083; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2085 = 10'h23 == ReadPtr[9:0] ? FifoCell_35 : _GEN_2084; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2086 = 10'h24 == ReadPtr[9:0] ? FifoCell_36 : _GEN_2085; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2087 = 10'h25 == ReadPtr[9:0] ? FifoCell_37 : _GEN_2086; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2088 = 10'h26 == ReadPtr[9:0] ? FifoCell_38 : _GEN_2087; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2089 = 10'h27 == ReadPtr[9:0] ? FifoCell_39 : _GEN_2088; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2090 = 10'h28 == ReadPtr[9:0] ? FifoCell_40 : _GEN_2089; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2091 = 10'h29 == ReadPtr[9:0] ? FifoCell_41 : _GEN_2090; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2092 = 10'h2a == ReadPtr[9:0] ? FifoCell_42 : _GEN_2091; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2093 = 10'h2b == ReadPtr[9:0] ? FifoCell_43 : _GEN_2092; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2094 = 10'h2c == ReadPtr[9:0] ? FifoCell_44 : _GEN_2093; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2095 = 10'h2d == ReadPtr[9:0] ? FifoCell_45 : _GEN_2094; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2096 = 10'h2e == ReadPtr[9:0] ? FifoCell_46 : _GEN_2095; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2097 = 10'h2f == ReadPtr[9:0] ? FifoCell_47 : _GEN_2096; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2098 = 10'h30 == ReadPtr[9:0] ? FifoCell_48 : _GEN_2097; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2099 = 10'h31 == ReadPtr[9:0] ? FifoCell_49 : _GEN_2098; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2100 = 10'h32 == ReadPtr[9:0] ? FifoCell_50 : _GEN_2099; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2101 = 10'h33 == ReadPtr[9:0] ? FifoCell_51 : _GEN_2100; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2102 = 10'h34 == ReadPtr[9:0] ? FifoCell_52 : _GEN_2101; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2103 = 10'h35 == ReadPtr[9:0] ? FifoCell_53 : _GEN_2102; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2104 = 10'h36 == ReadPtr[9:0] ? FifoCell_54 : _GEN_2103; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2105 = 10'h37 == ReadPtr[9:0] ? FifoCell_55 : _GEN_2104; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2106 = 10'h38 == ReadPtr[9:0] ? FifoCell_56 : _GEN_2105; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2107 = 10'h39 == ReadPtr[9:0] ? FifoCell_57 : _GEN_2106; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2108 = 10'h3a == ReadPtr[9:0] ? FifoCell_58 : _GEN_2107; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2109 = 10'h3b == ReadPtr[9:0] ? FifoCell_59 : _GEN_2108; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2110 = 10'h3c == ReadPtr[9:0] ? FifoCell_60 : _GEN_2109; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2111 = 10'h3d == ReadPtr[9:0] ? FifoCell_61 : _GEN_2110; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2112 = 10'h3e == ReadPtr[9:0] ? FifoCell_62 : _GEN_2111; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2113 = 10'h3f == ReadPtr[9:0] ? FifoCell_63 : _GEN_2112; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2114 = 10'h40 == ReadPtr[9:0] ? FifoCell_64 : _GEN_2113; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2115 = 10'h41 == ReadPtr[9:0] ? FifoCell_65 : _GEN_2114; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2116 = 10'h42 == ReadPtr[9:0] ? FifoCell_66 : _GEN_2115; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2117 = 10'h43 == ReadPtr[9:0] ? FifoCell_67 : _GEN_2116; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2118 = 10'h44 == ReadPtr[9:0] ? FifoCell_68 : _GEN_2117; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2119 = 10'h45 == ReadPtr[9:0] ? FifoCell_69 : _GEN_2118; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2120 = 10'h46 == ReadPtr[9:0] ? FifoCell_70 : _GEN_2119; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2121 = 10'h47 == ReadPtr[9:0] ? FifoCell_71 : _GEN_2120; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2122 = 10'h48 == ReadPtr[9:0] ? FifoCell_72 : _GEN_2121; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2123 = 10'h49 == ReadPtr[9:0] ? FifoCell_73 : _GEN_2122; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2124 = 10'h4a == ReadPtr[9:0] ? FifoCell_74 : _GEN_2123; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2125 = 10'h4b == ReadPtr[9:0] ? FifoCell_75 : _GEN_2124; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2126 = 10'h4c == ReadPtr[9:0] ? FifoCell_76 : _GEN_2125; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2127 = 10'h4d == ReadPtr[9:0] ? FifoCell_77 : _GEN_2126; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2128 = 10'h4e == ReadPtr[9:0] ? FifoCell_78 : _GEN_2127; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2129 = 10'h4f == ReadPtr[9:0] ? FifoCell_79 : _GEN_2128; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2130 = 10'h50 == ReadPtr[9:0] ? FifoCell_80 : _GEN_2129; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2131 = 10'h51 == ReadPtr[9:0] ? FifoCell_81 : _GEN_2130; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2132 = 10'h52 == ReadPtr[9:0] ? FifoCell_82 : _GEN_2131; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2133 = 10'h53 == ReadPtr[9:0] ? FifoCell_83 : _GEN_2132; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2134 = 10'h54 == ReadPtr[9:0] ? FifoCell_84 : _GEN_2133; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2135 = 10'h55 == ReadPtr[9:0] ? FifoCell_85 : _GEN_2134; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2136 = 10'h56 == ReadPtr[9:0] ? FifoCell_86 : _GEN_2135; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2137 = 10'h57 == ReadPtr[9:0] ? FifoCell_87 : _GEN_2136; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2138 = 10'h58 == ReadPtr[9:0] ? FifoCell_88 : _GEN_2137; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2139 = 10'h59 == ReadPtr[9:0] ? FifoCell_89 : _GEN_2138; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2140 = 10'h5a == ReadPtr[9:0] ? FifoCell_90 : _GEN_2139; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2141 = 10'h5b == ReadPtr[9:0] ? FifoCell_91 : _GEN_2140; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2142 = 10'h5c == ReadPtr[9:0] ? FifoCell_92 : _GEN_2141; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2143 = 10'h5d == ReadPtr[9:0] ? FifoCell_93 : _GEN_2142; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2144 = 10'h5e == ReadPtr[9:0] ? FifoCell_94 : _GEN_2143; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2145 = 10'h5f == ReadPtr[9:0] ? FifoCell_95 : _GEN_2144; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2146 = 10'h60 == ReadPtr[9:0] ? FifoCell_96 : _GEN_2145; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2147 = 10'h61 == ReadPtr[9:0] ? FifoCell_97 : _GEN_2146; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2148 = 10'h62 == ReadPtr[9:0] ? FifoCell_98 : _GEN_2147; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2149 = 10'h63 == ReadPtr[9:0] ? FifoCell_99 : _GEN_2148; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2150 = 10'h64 == ReadPtr[9:0] ? FifoCell_100 : _GEN_2149; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2151 = 10'h65 == ReadPtr[9:0] ? FifoCell_101 : _GEN_2150; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2152 = 10'h66 == ReadPtr[9:0] ? FifoCell_102 : _GEN_2151; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2153 = 10'h67 == ReadPtr[9:0] ? FifoCell_103 : _GEN_2152; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2154 = 10'h68 == ReadPtr[9:0] ? FifoCell_104 : _GEN_2153; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2155 = 10'h69 == ReadPtr[9:0] ? FifoCell_105 : _GEN_2154; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2156 = 10'h6a == ReadPtr[9:0] ? FifoCell_106 : _GEN_2155; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2157 = 10'h6b == ReadPtr[9:0] ? FifoCell_107 : _GEN_2156; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2158 = 10'h6c == ReadPtr[9:0] ? FifoCell_108 : _GEN_2157; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2159 = 10'h6d == ReadPtr[9:0] ? FifoCell_109 : _GEN_2158; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2160 = 10'h6e == ReadPtr[9:0] ? FifoCell_110 : _GEN_2159; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2161 = 10'h6f == ReadPtr[9:0] ? FifoCell_111 : _GEN_2160; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2162 = 10'h70 == ReadPtr[9:0] ? FifoCell_112 : _GEN_2161; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2163 = 10'h71 == ReadPtr[9:0] ? FifoCell_113 : _GEN_2162; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2164 = 10'h72 == ReadPtr[9:0] ? FifoCell_114 : _GEN_2163; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2165 = 10'h73 == ReadPtr[9:0] ? FifoCell_115 : _GEN_2164; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2166 = 10'h74 == ReadPtr[9:0] ? FifoCell_116 : _GEN_2165; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2167 = 10'h75 == ReadPtr[9:0] ? FifoCell_117 : _GEN_2166; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2168 = 10'h76 == ReadPtr[9:0] ? FifoCell_118 : _GEN_2167; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2169 = 10'h77 == ReadPtr[9:0] ? FifoCell_119 : _GEN_2168; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2170 = 10'h78 == ReadPtr[9:0] ? FifoCell_120 : _GEN_2169; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2171 = 10'h79 == ReadPtr[9:0] ? FifoCell_121 : _GEN_2170; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2172 = 10'h7a == ReadPtr[9:0] ? FifoCell_122 : _GEN_2171; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2173 = 10'h7b == ReadPtr[9:0] ? FifoCell_123 : _GEN_2172; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2174 = 10'h7c == ReadPtr[9:0] ? FifoCell_124 : _GEN_2173; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2175 = 10'h7d == ReadPtr[9:0] ? FifoCell_125 : _GEN_2174; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2176 = 10'h7e == ReadPtr[9:0] ? FifoCell_126 : _GEN_2175; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2177 = 10'h7f == ReadPtr[9:0] ? FifoCell_127 : _GEN_2176; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2178 = 10'h80 == ReadPtr[9:0] ? FifoCell_128 : _GEN_2177; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2179 = 10'h81 == ReadPtr[9:0] ? FifoCell_129 : _GEN_2178; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2180 = 10'h82 == ReadPtr[9:0] ? FifoCell_130 : _GEN_2179; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2181 = 10'h83 == ReadPtr[9:0] ? FifoCell_131 : _GEN_2180; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2182 = 10'h84 == ReadPtr[9:0] ? FifoCell_132 : _GEN_2181; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2183 = 10'h85 == ReadPtr[9:0] ? FifoCell_133 : _GEN_2182; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2184 = 10'h86 == ReadPtr[9:0] ? FifoCell_134 : _GEN_2183; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2185 = 10'h87 == ReadPtr[9:0] ? FifoCell_135 : _GEN_2184; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2186 = 10'h88 == ReadPtr[9:0] ? FifoCell_136 : _GEN_2185; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2187 = 10'h89 == ReadPtr[9:0] ? FifoCell_137 : _GEN_2186; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2188 = 10'h8a == ReadPtr[9:0] ? FifoCell_138 : _GEN_2187; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2189 = 10'h8b == ReadPtr[9:0] ? FifoCell_139 : _GEN_2188; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2190 = 10'h8c == ReadPtr[9:0] ? FifoCell_140 : _GEN_2189; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2191 = 10'h8d == ReadPtr[9:0] ? FifoCell_141 : _GEN_2190; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2192 = 10'h8e == ReadPtr[9:0] ? FifoCell_142 : _GEN_2191; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2193 = 10'h8f == ReadPtr[9:0] ? FifoCell_143 : _GEN_2192; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2194 = 10'h90 == ReadPtr[9:0] ? FifoCell_144 : _GEN_2193; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2195 = 10'h91 == ReadPtr[9:0] ? FifoCell_145 : _GEN_2194; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2196 = 10'h92 == ReadPtr[9:0] ? FifoCell_146 : _GEN_2195; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2197 = 10'h93 == ReadPtr[9:0] ? FifoCell_147 : _GEN_2196; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2198 = 10'h94 == ReadPtr[9:0] ? FifoCell_148 : _GEN_2197; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2199 = 10'h95 == ReadPtr[9:0] ? FifoCell_149 : _GEN_2198; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2200 = 10'h96 == ReadPtr[9:0] ? FifoCell_150 : _GEN_2199; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2201 = 10'h97 == ReadPtr[9:0] ? FifoCell_151 : _GEN_2200; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2202 = 10'h98 == ReadPtr[9:0] ? FifoCell_152 : _GEN_2201; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2203 = 10'h99 == ReadPtr[9:0] ? FifoCell_153 : _GEN_2202; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2204 = 10'h9a == ReadPtr[9:0] ? FifoCell_154 : _GEN_2203; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2205 = 10'h9b == ReadPtr[9:0] ? FifoCell_155 : _GEN_2204; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2206 = 10'h9c == ReadPtr[9:0] ? FifoCell_156 : _GEN_2205; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2207 = 10'h9d == ReadPtr[9:0] ? FifoCell_157 : _GEN_2206; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2208 = 10'h9e == ReadPtr[9:0] ? FifoCell_158 : _GEN_2207; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2209 = 10'h9f == ReadPtr[9:0] ? FifoCell_159 : _GEN_2208; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2210 = 10'ha0 == ReadPtr[9:0] ? FifoCell_160 : _GEN_2209; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2211 = 10'ha1 == ReadPtr[9:0] ? FifoCell_161 : _GEN_2210; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2212 = 10'ha2 == ReadPtr[9:0] ? FifoCell_162 : _GEN_2211; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2213 = 10'ha3 == ReadPtr[9:0] ? FifoCell_163 : _GEN_2212; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2214 = 10'ha4 == ReadPtr[9:0] ? FifoCell_164 : _GEN_2213; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2215 = 10'ha5 == ReadPtr[9:0] ? FifoCell_165 : _GEN_2214; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2216 = 10'ha6 == ReadPtr[9:0] ? FifoCell_166 : _GEN_2215; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2217 = 10'ha7 == ReadPtr[9:0] ? FifoCell_167 : _GEN_2216; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2218 = 10'ha8 == ReadPtr[9:0] ? FifoCell_168 : _GEN_2217; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2219 = 10'ha9 == ReadPtr[9:0] ? FifoCell_169 : _GEN_2218; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2220 = 10'haa == ReadPtr[9:0] ? FifoCell_170 : _GEN_2219; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2221 = 10'hab == ReadPtr[9:0] ? FifoCell_171 : _GEN_2220; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2222 = 10'hac == ReadPtr[9:0] ? FifoCell_172 : _GEN_2221; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2223 = 10'had == ReadPtr[9:0] ? FifoCell_173 : _GEN_2222; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2224 = 10'hae == ReadPtr[9:0] ? FifoCell_174 : _GEN_2223; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2225 = 10'haf == ReadPtr[9:0] ? FifoCell_175 : _GEN_2224; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2226 = 10'hb0 == ReadPtr[9:0] ? FifoCell_176 : _GEN_2225; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2227 = 10'hb1 == ReadPtr[9:0] ? FifoCell_177 : _GEN_2226; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2228 = 10'hb2 == ReadPtr[9:0] ? FifoCell_178 : _GEN_2227; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2229 = 10'hb3 == ReadPtr[9:0] ? FifoCell_179 : _GEN_2228; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2230 = 10'hb4 == ReadPtr[9:0] ? FifoCell_180 : _GEN_2229; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2231 = 10'hb5 == ReadPtr[9:0] ? FifoCell_181 : _GEN_2230; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2232 = 10'hb6 == ReadPtr[9:0] ? FifoCell_182 : _GEN_2231; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2233 = 10'hb7 == ReadPtr[9:0] ? FifoCell_183 : _GEN_2232; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2234 = 10'hb8 == ReadPtr[9:0] ? FifoCell_184 : _GEN_2233; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2235 = 10'hb9 == ReadPtr[9:0] ? FifoCell_185 : _GEN_2234; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2236 = 10'hba == ReadPtr[9:0] ? FifoCell_186 : _GEN_2235; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2237 = 10'hbb == ReadPtr[9:0] ? FifoCell_187 : _GEN_2236; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2238 = 10'hbc == ReadPtr[9:0] ? FifoCell_188 : _GEN_2237; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2239 = 10'hbd == ReadPtr[9:0] ? FifoCell_189 : _GEN_2238; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2240 = 10'hbe == ReadPtr[9:0] ? FifoCell_190 : _GEN_2239; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2241 = 10'hbf == ReadPtr[9:0] ? FifoCell_191 : _GEN_2240; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2242 = 10'hc0 == ReadPtr[9:0] ? FifoCell_192 : _GEN_2241; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2243 = 10'hc1 == ReadPtr[9:0] ? FifoCell_193 : _GEN_2242; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2244 = 10'hc2 == ReadPtr[9:0] ? FifoCell_194 : _GEN_2243; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2245 = 10'hc3 == ReadPtr[9:0] ? FifoCell_195 : _GEN_2244; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2246 = 10'hc4 == ReadPtr[9:0] ? FifoCell_196 : _GEN_2245; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2247 = 10'hc5 == ReadPtr[9:0] ? FifoCell_197 : _GEN_2246; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2248 = 10'hc6 == ReadPtr[9:0] ? FifoCell_198 : _GEN_2247; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2249 = 10'hc7 == ReadPtr[9:0] ? FifoCell_199 : _GEN_2248; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2250 = 10'hc8 == ReadPtr[9:0] ? FifoCell_200 : _GEN_2249; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2251 = 10'hc9 == ReadPtr[9:0] ? FifoCell_201 : _GEN_2250; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2252 = 10'hca == ReadPtr[9:0] ? FifoCell_202 : _GEN_2251; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2253 = 10'hcb == ReadPtr[9:0] ? FifoCell_203 : _GEN_2252; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2254 = 10'hcc == ReadPtr[9:0] ? FifoCell_204 : _GEN_2253; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2255 = 10'hcd == ReadPtr[9:0] ? FifoCell_205 : _GEN_2254; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2256 = 10'hce == ReadPtr[9:0] ? FifoCell_206 : _GEN_2255; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2257 = 10'hcf == ReadPtr[9:0] ? FifoCell_207 : _GEN_2256; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2258 = 10'hd0 == ReadPtr[9:0] ? FifoCell_208 : _GEN_2257; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2259 = 10'hd1 == ReadPtr[9:0] ? FifoCell_209 : _GEN_2258; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2260 = 10'hd2 == ReadPtr[9:0] ? FifoCell_210 : _GEN_2259; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2261 = 10'hd3 == ReadPtr[9:0] ? FifoCell_211 : _GEN_2260; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2262 = 10'hd4 == ReadPtr[9:0] ? FifoCell_212 : _GEN_2261; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2263 = 10'hd5 == ReadPtr[9:0] ? FifoCell_213 : _GEN_2262; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2264 = 10'hd6 == ReadPtr[9:0] ? FifoCell_214 : _GEN_2263; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2265 = 10'hd7 == ReadPtr[9:0] ? FifoCell_215 : _GEN_2264; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2266 = 10'hd8 == ReadPtr[9:0] ? FifoCell_216 : _GEN_2265; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2267 = 10'hd9 == ReadPtr[9:0] ? FifoCell_217 : _GEN_2266; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2268 = 10'hda == ReadPtr[9:0] ? FifoCell_218 : _GEN_2267; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2269 = 10'hdb == ReadPtr[9:0] ? FifoCell_219 : _GEN_2268; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2270 = 10'hdc == ReadPtr[9:0] ? FifoCell_220 : _GEN_2269; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2271 = 10'hdd == ReadPtr[9:0] ? FifoCell_221 : _GEN_2270; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2272 = 10'hde == ReadPtr[9:0] ? FifoCell_222 : _GEN_2271; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2273 = 10'hdf == ReadPtr[9:0] ? FifoCell_223 : _GEN_2272; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2274 = 10'he0 == ReadPtr[9:0] ? FifoCell_224 : _GEN_2273; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2275 = 10'he1 == ReadPtr[9:0] ? FifoCell_225 : _GEN_2274; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2276 = 10'he2 == ReadPtr[9:0] ? FifoCell_226 : _GEN_2275; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2277 = 10'he3 == ReadPtr[9:0] ? FifoCell_227 : _GEN_2276; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2278 = 10'he4 == ReadPtr[9:0] ? FifoCell_228 : _GEN_2277; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2279 = 10'he5 == ReadPtr[9:0] ? FifoCell_229 : _GEN_2278; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2280 = 10'he6 == ReadPtr[9:0] ? FifoCell_230 : _GEN_2279; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2281 = 10'he7 == ReadPtr[9:0] ? FifoCell_231 : _GEN_2280; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2282 = 10'he8 == ReadPtr[9:0] ? FifoCell_232 : _GEN_2281; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2283 = 10'he9 == ReadPtr[9:0] ? FifoCell_233 : _GEN_2282; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2284 = 10'hea == ReadPtr[9:0] ? FifoCell_234 : _GEN_2283; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2285 = 10'heb == ReadPtr[9:0] ? FifoCell_235 : _GEN_2284; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2286 = 10'hec == ReadPtr[9:0] ? FifoCell_236 : _GEN_2285; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2287 = 10'hed == ReadPtr[9:0] ? FifoCell_237 : _GEN_2286; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2288 = 10'hee == ReadPtr[9:0] ? FifoCell_238 : _GEN_2287; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2289 = 10'hef == ReadPtr[9:0] ? FifoCell_239 : _GEN_2288; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2290 = 10'hf0 == ReadPtr[9:0] ? FifoCell_240 : _GEN_2289; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2291 = 10'hf1 == ReadPtr[9:0] ? FifoCell_241 : _GEN_2290; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2292 = 10'hf2 == ReadPtr[9:0] ? FifoCell_242 : _GEN_2291; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2293 = 10'hf3 == ReadPtr[9:0] ? FifoCell_243 : _GEN_2292; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2294 = 10'hf4 == ReadPtr[9:0] ? FifoCell_244 : _GEN_2293; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2295 = 10'hf5 == ReadPtr[9:0] ? FifoCell_245 : _GEN_2294; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2296 = 10'hf6 == ReadPtr[9:0] ? FifoCell_246 : _GEN_2295; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2297 = 10'hf7 == ReadPtr[9:0] ? FifoCell_247 : _GEN_2296; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2298 = 10'hf8 == ReadPtr[9:0] ? FifoCell_248 : _GEN_2297; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2299 = 10'hf9 == ReadPtr[9:0] ? FifoCell_249 : _GEN_2298; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2300 = 10'hfa == ReadPtr[9:0] ? FifoCell_250 : _GEN_2299; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2301 = 10'hfb == ReadPtr[9:0] ? FifoCell_251 : _GEN_2300; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2302 = 10'hfc == ReadPtr[9:0] ? FifoCell_252 : _GEN_2301; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2303 = 10'hfd == ReadPtr[9:0] ? FifoCell_253 : _GEN_2302; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2304 = 10'hfe == ReadPtr[9:0] ? FifoCell_254 : _GEN_2303; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2305 = 10'hff == ReadPtr[9:0] ? FifoCell_255 : _GEN_2304; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2306 = 10'h100 == ReadPtr[9:0] ? FifoCell_256 : _GEN_2305; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2307 = 10'h101 == ReadPtr[9:0] ? FifoCell_257 : _GEN_2306; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2308 = 10'h102 == ReadPtr[9:0] ? FifoCell_258 : _GEN_2307; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2309 = 10'h103 == ReadPtr[9:0] ? FifoCell_259 : _GEN_2308; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2310 = 10'h104 == ReadPtr[9:0] ? FifoCell_260 : _GEN_2309; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2311 = 10'h105 == ReadPtr[9:0] ? FifoCell_261 : _GEN_2310; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2312 = 10'h106 == ReadPtr[9:0] ? FifoCell_262 : _GEN_2311; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2313 = 10'h107 == ReadPtr[9:0] ? FifoCell_263 : _GEN_2312; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2314 = 10'h108 == ReadPtr[9:0] ? FifoCell_264 : _GEN_2313; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2315 = 10'h109 == ReadPtr[9:0] ? FifoCell_265 : _GEN_2314; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2316 = 10'h10a == ReadPtr[9:0] ? FifoCell_266 : _GEN_2315; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2317 = 10'h10b == ReadPtr[9:0] ? FifoCell_267 : _GEN_2316; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2318 = 10'h10c == ReadPtr[9:0] ? FifoCell_268 : _GEN_2317; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2319 = 10'h10d == ReadPtr[9:0] ? FifoCell_269 : _GEN_2318; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2320 = 10'h10e == ReadPtr[9:0] ? FifoCell_270 : _GEN_2319; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2321 = 10'h10f == ReadPtr[9:0] ? FifoCell_271 : _GEN_2320; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2322 = 10'h110 == ReadPtr[9:0] ? FifoCell_272 : _GEN_2321; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2323 = 10'h111 == ReadPtr[9:0] ? FifoCell_273 : _GEN_2322; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2324 = 10'h112 == ReadPtr[9:0] ? FifoCell_274 : _GEN_2323; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2325 = 10'h113 == ReadPtr[9:0] ? FifoCell_275 : _GEN_2324; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2326 = 10'h114 == ReadPtr[9:0] ? FifoCell_276 : _GEN_2325; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2327 = 10'h115 == ReadPtr[9:0] ? FifoCell_277 : _GEN_2326; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2328 = 10'h116 == ReadPtr[9:0] ? FifoCell_278 : _GEN_2327; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2329 = 10'h117 == ReadPtr[9:0] ? FifoCell_279 : _GEN_2328; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2330 = 10'h118 == ReadPtr[9:0] ? FifoCell_280 : _GEN_2329; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2331 = 10'h119 == ReadPtr[9:0] ? FifoCell_281 : _GEN_2330; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2332 = 10'h11a == ReadPtr[9:0] ? FifoCell_282 : _GEN_2331; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2333 = 10'h11b == ReadPtr[9:0] ? FifoCell_283 : _GEN_2332; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2334 = 10'h11c == ReadPtr[9:0] ? FifoCell_284 : _GEN_2333; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2335 = 10'h11d == ReadPtr[9:0] ? FifoCell_285 : _GEN_2334; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2336 = 10'h11e == ReadPtr[9:0] ? FifoCell_286 : _GEN_2335; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2337 = 10'h11f == ReadPtr[9:0] ? FifoCell_287 : _GEN_2336; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2338 = 10'h120 == ReadPtr[9:0] ? FifoCell_288 : _GEN_2337; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2339 = 10'h121 == ReadPtr[9:0] ? FifoCell_289 : _GEN_2338; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2340 = 10'h122 == ReadPtr[9:0] ? FifoCell_290 : _GEN_2339; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2341 = 10'h123 == ReadPtr[9:0] ? FifoCell_291 : _GEN_2340; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2342 = 10'h124 == ReadPtr[9:0] ? FifoCell_292 : _GEN_2341; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2343 = 10'h125 == ReadPtr[9:0] ? FifoCell_293 : _GEN_2342; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2344 = 10'h126 == ReadPtr[9:0] ? FifoCell_294 : _GEN_2343; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2345 = 10'h127 == ReadPtr[9:0] ? FifoCell_295 : _GEN_2344; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2346 = 10'h128 == ReadPtr[9:0] ? FifoCell_296 : _GEN_2345; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2347 = 10'h129 == ReadPtr[9:0] ? FifoCell_297 : _GEN_2346; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2348 = 10'h12a == ReadPtr[9:0] ? FifoCell_298 : _GEN_2347; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2349 = 10'h12b == ReadPtr[9:0] ? FifoCell_299 : _GEN_2348; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2350 = 10'h12c == ReadPtr[9:0] ? FifoCell_300 : _GEN_2349; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2351 = 10'h12d == ReadPtr[9:0] ? FifoCell_301 : _GEN_2350; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2352 = 10'h12e == ReadPtr[9:0] ? FifoCell_302 : _GEN_2351; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2353 = 10'h12f == ReadPtr[9:0] ? FifoCell_303 : _GEN_2352; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2354 = 10'h130 == ReadPtr[9:0] ? FifoCell_304 : _GEN_2353; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2355 = 10'h131 == ReadPtr[9:0] ? FifoCell_305 : _GEN_2354; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2356 = 10'h132 == ReadPtr[9:0] ? FifoCell_306 : _GEN_2355; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2357 = 10'h133 == ReadPtr[9:0] ? FifoCell_307 : _GEN_2356; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2358 = 10'h134 == ReadPtr[9:0] ? FifoCell_308 : _GEN_2357; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2359 = 10'h135 == ReadPtr[9:0] ? FifoCell_309 : _GEN_2358; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2360 = 10'h136 == ReadPtr[9:0] ? FifoCell_310 : _GEN_2359; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2361 = 10'h137 == ReadPtr[9:0] ? FifoCell_311 : _GEN_2360; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2362 = 10'h138 == ReadPtr[9:0] ? FifoCell_312 : _GEN_2361; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2363 = 10'h139 == ReadPtr[9:0] ? FifoCell_313 : _GEN_2362; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2364 = 10'h13a == ReadPtr[9:0] ? FifoCell_314 : _GEN_2363; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2365 = 10'h13b == ReadPtr[9:0] ? FifoCell_315 : _GEN_2364; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2366 = 10'h13c == ReadPtr[9:0] ? FifoCell_316 : _GEN_2365; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2367 = 10'h13d == ReadPtr[9:0] ? FifoCell_317 : _GEN_2366; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2368 = 10'h13e == ReadPtr[9:0] ? FifoCell_318 : _GEN_2367; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2369 = 10'h13f == ReadPtr[9:0] ? FifoCell_319 : _GEN_2368; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2370 = 10'h140 == ReadPtr[9:0] ? FifoCell_320 : _GEN_2369; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2371 = 10'h141 == ReadPtr[9:0] ? FifoCell_321 : _GEN_2370; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2372 = 10'h142 == ReadPtr[9:0] ? FifoCell_322 : _GEN_2371; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2373 = 10'h143 == ReadPtr[9:0] ? FifoCell_323 : _GEN_2372; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2374 = 10'h144 == ReadPtr[9:0] ? FifoCell_324 : _GEN_2373; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2375 = 10'h145 == ReadPtr[9:0] ? FifoCell_325 : _GEN_2374; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2376 = 10'h146 == ReadPtr[9:0] ? FifoCell_326 : _GEN_2375; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2377 = 10'h147 == ReadPtr[9:0] ? FifoCell_327 : _GEN_2376; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2378 = 10'h148 == ReadPtr[9:0] ? FifoCell_328 : _GEN_2377; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2379 = 10'h149 == ReadPtr[9:0] ? FifoCell_329 : _GEN_2378; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2380 = 10'h14a == ReadPtr[9:0] ? FifoCell_330 : _GEN_2379; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2381 = 10'h14b == ReadPtr[9:0] ? FifoCell_331 : _GEN_2380; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2382 = 10'h14c == ReadPtr[9:0] ? FifoCell_332 : _GEN_2381; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2383 = 10'h14d == ReadPtr[9:0] ? FifoCell_333 : _GEN_2382; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2384 = 10'h14e == ReadPtr[9:0] ? FifoCell_334 : _GEN_2383; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2385 = 10'h14f == ReadPtr[9:0] ? FifoCell_335 : _GEN_2384; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2386 = 10'h150 == ReadPtr[9:0] ? FifoCell_336 : _GEN_2385; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2387 = 10'h151 == ReadPtr[9:0] ? FifoCell_337 : _GEN_2386; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2388 = 10'h152 == ReadPtr[9:0] ? FifoCell_338 : _GEN_2387; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2389 = 10'h153 == ReadPtr[9:0] ? FifoCell_339 : _GEN_2388; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2390 = 10'h154 == ReadPtr[9:0] ? FifoCell_340 : _GEN_2389; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2391 = 10'h155 == ReadPtr[9:0] ? FifoCell_341 : _GEN_2390; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2392 = 10'h156 == ReadPtr[9:0] ? FifoCell_342 : _GEN_2391; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2393 = 10'h157 == ReadPtr[9:0] ? FifoCell_343 : _GEN_2392; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2394 = 10'h158 == ReadPtr[9:0] ? FifoCell_344 : _GEN_2393; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2395 = 10'h159 == ReadPtr[9:0] ? FifoCell_345 : _GEN_2394; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2396 = 10'h15a == ReadPtr[9:0] ? FifoCell_346 : _GEN_2395; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2397 = 10'h15b == ReadPtr[9:0] ? FifoCell_347 : _GEN_2396; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2398 = 10'h15c == ReadPtr[9:0] ? FifoCell_348 : _GEN_2397; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2399 = 10'h15d == ReadPtr[9:0] ? FifoCell_349 : _GEN_2398; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2400 = 10'h15e == ReadPtr[9:0] ? FifoCell_350 : _GEN_2399; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2401 = 10'h15f == ReadPtr[9:0] ? FifoCell_351 : _GEN_2400; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2402 = 10'h160 == ReadPtr[9:0] ? FifoCell_352 : _GEN_2401; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2403 = 10'h161 == ReadPtr[9:0] ? FifoCell_353 : _GEN_2402; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2404 = 10'h162 == ReadPtr[9:0] ? FifoCell_354 : _GEN_2403; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2405 = 10'h163 == ReadPtr[9:0] ? FifoCell_355 : _GEN_2404; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2406 = 10'h164 == ReadPtr[9:0] ? FifoCell_356 : _GEN_2405; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2407 = 10'h165 == ReadPtr[9:0] ? FifoCell_357 : _GEN_2406; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2408 = 10'h166 == ReadPtr[9:0] ? FifoCell_358 : _GEN_2407; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2409 = 10'h167 == ReadPtr[9:0] ? FifoCell_359 : _GEN_2408; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2410 = 10'h168 == ReadPtr[9:0] ? FifoCell_360 : _GEN_2409; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2411 = 10'h169 == ReadPtr[9:0] ? FifoCell_361 : _GEN_2410; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2412 = 10'h16a == ReadPtr[9:0] ? FifoCell_362 : _GEN_2411; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2413 = 10'h16b == ReadPtr[9:0] ? FifoCell_363 : _GEN_2412; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2414 = 10'h16c == ReadPtr[9:0] ? FifoCell_364 : _GEN_2413; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2415 = 10'h16d == ReadPtr[9:0] ? FifoCell_365 : _GEN_2414; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2416 = 10'h16e == ReadPtr[9:0] ? FifoCell_366 : _GEN_2415; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2417 = 10'h16f == ReadPtr[9:0] ? FifoCell_367 : _GEN_2416; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2418 = 10'h170 == ReadPtr[9:0] ? FifoCell_368 : _GEN_2417; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2419 = 10'h171 == ReadPtr[9:0] ? FifoCell_369 : _GEN_2418; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2420 = 10'h172 == ReadPtr[9:0] ? FifoCell_370 : _GEN_2419; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2421 = 10'h173 == ReadPtr[9:0] ? FifoCell_371 : _GEN_2420; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2422 = 10'h174 == ReadPtr[9:0] ? FifoCell_372 : _GEN_2421; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2423 = 10'h175 == ReadPtr[9:0] ? FifoCell_373 : _GEN_2422; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2424 = 10'h176 == ReadPtr[9:0] ? FifoCell_374 : _GEN_2423; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2425 = 10'h177 == ReadPtr[9:0] ? FifoCell_375 : _GEN_2424; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2426 = 10'h178 == ReadPtr[9:0] ? FifoCell_376 : _GEN_2425; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2427 = 10'h179 == ReadPtr[9:0] ? FifoCell_377 : _GEN_2426; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2428 = 10'h17a == ReadPtr[9:0] ? FifoCell_378 : _GEN_2427; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2429 = 10'h17b == ReadPtr[9:0] ? FifoCell_379 : _GEN_2428; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2430 = 10'h17c == ReadPtr[9:0] ? FifoCell_380 : _GEN_2429; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2431 = 10'h17d == ReadPtr[9:0] ? FifoCell_381 : _GEN_2430; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2432 = 10'h17e == ReadPtr[9:0] ? FifoCell_382 : _GEN_2431; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2433 = 10'h17f == ReadPtr[9:0] ? FifoCell_383 : _GEN_2432; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2434 = 10'h180 == ReadPtr[9:0] ? FifoCell_384 : _GEN_2433; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2435 = 10'h181 == ReadPtr[9:0] ? FifoCell_385 : _GEN_2434; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2436 = 10'h182 == ReadPtr[9:0] ? FifoCell_386 : _GEN_2435; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2437 = 10'h183 == ReadPtr[9:0] ? FifoCell_387 : _GEN_2436; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2438 = 10'h184 == ReadPtr[9:0] ? FifoCell_388 : _GEN_2437; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2439 = 10'h185 == ReadPtr[9:0] ? FifoCell_389 : _GEN_2438; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2440 = 10'h186 == ReadPtr[9:0] ? FifoCell_390 : _GEN_2439; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2441 = 10'h187 == ReadPtr[9:0] ? FifoCell_391 : _GEN_2440; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2442 = 10'h188 == ReadPtr[9:0] ? FifoCell_392 : _GEN_2441; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2443 = 10'h189 == ReadPtr[9:0] ? FifoCell_393 : _GEN_2442; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2444 = 10'h18a == ReadPtr[9:0] ? FifoCell_394 : _GEN_2443; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2445 = 10'h18b == ReadPtr[9:0] ? FifoCell_395 : _GEN_2444; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2446 = 10'h18c == ReadPtr[9:0] ? FifoCell_396 : _GEN_2445; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2447 = 10'h18d == ReadPtr[9:0] ? FifoCell_397 : _GEN_2446; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2448 = 10'h18e == ReadPtr[9:0] ? FifoCell_398 : _GEN_2447; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2449 = 10'h18f == ReadPtr[9:0] ? FifoCell_399 : _GEN_2448; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2450 = 10'h190 == ReadPtr[9:0] ? FifoCell_400 : _GEN_2449; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2451 = 10'h191 == ReadPtr[9:0] ? FifoCell_401 : _GEN_2450; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2452 = 10'h192 == ReadPtr[9:0] ? FifoCell_402 : _GEN_2451; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2453 = 10'h193 == ReadPtr[9:0] ? FifoCell_403 : _GEN_2452; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2454 = 10'h194 == ReadPtr[9:0] ? FifoCell_404 : _GEN_2453; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2455 = 10'h195 == ReadPtr[9:0] ? FifoCell_405 : _GEN_2454; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2456 = 10'h196 == ReadPtr[9:0] ? FifoCell_406 : _GEN_2455; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2457 = 10'h197 == ReadPtr[9:0] ? FifoCell_407 : _GEN_2456; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2458 = 10'h198 == ReadPtr[9:0] ? FifoCell_408 : _GEN_2457; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2459 = 10'h199 == ReadPtr[9:0] ? FifoCell_409 : _GEN_2458; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2460 = 10'h19a == ReadPtr[9:0] ? FifoCell_410 : _GEN_2459; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2461 = 10'h19b == ReadPtr[9:0] ? FifoCell_411 : _GEN_2460; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2462 = 10'h19c == ReadPtr[9:0] ? FifoCell_412 : _GEN_2461; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2463 = 10'h19d == ReadPtr[9:0] ? FifoCell_413 : _GEN_2462; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2464 = 10'h19e == ReadPtr[9:0] ? FifoCell_414 : _GEN_2463; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2465 = 10'h19f == ReadPtr[9:0] ? FifoCell_415 : _GEN_2464; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2466 = 10'h1a0 == ReadPtr[9:0] ? FifoCell_416 : _GEN_2465; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2467 = 10'h1a1 == ReadPtr[9:0] ? FifoCell_417 : _GEN_2466; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2468 = 10'h1a2 == ReadPtr[9:0] ? FifoCell_418 : _GEN_2467; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2469 = 10'h1a3 == ReadPtr[9:0] ? FifoCell_419 : _GEN_2468; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2470 = 10'h1a4 == ReadPtr[9:0] ? FifoCell_420 : _GEN_2469; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2471 = 10'h1a5 == ReadPtr[9:0] ? FifoCell_421 : _GEN_2470; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2472 = 10'h1a6 == ReadPtr[9:0] ? FifoCell_422 : _GEN_2471; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2473 = 10'h1a7 == ReadPtr[9:0] ? FifoCell_423 : _GEN_2472; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2474 = 10'h1a8 == ReadPtr[9:0] ? FifoCell_424 : _GEN_2473; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2475 = 10'h1a9 == ReadPtr[9:0] ? FifoCell_425 : _GEN_2474; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2476 = 10'h1aa == ReadPtr[9:0] ? FifoCell_426 : _GEN_2475; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2477 = 10'h1ab == ReadPtr[9:0] ? FifoCell_427 : _GEN_2476; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2478 = 10'h1ac == ReadPtr[9:0] ? FifoCell_428 : _GEN_2477; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2479 = 10'h1ad == ReadPtr[9:0] ? FifoCell_429 : _GEN_2478; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2480 = 10'h1ae == ReadPtr[9:0] ? FifoCell_430 : _GEN_2479; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2481 = 10'h1af == ReadPtr[9:0] ? FifoCell_431 : _GEN_2480; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2482 = 10'h1b0 == ReadPtr[9:0] ? FifoCell_432 : _GEN_2481; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2483 = 10'h1b1 == ReadPtr[9:0] ? FifoCell_433 : _GEN_2482; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2484 = 10'h1b2 == ReadPtr[9:0] ? FifoCell_434 : _GEN_2483; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2485 = 10'h1b3 == ReadPtr[9:0] ? FifoCell_435 : _GEN_2484; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2486 = 10'h1b4 == ReadPtr[9:0] ? FifoCell_436 : _GEN_2485; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2487 = 10'h1b5 == ReadPtr[9:0] ? FifoCell_437 : _GEN_2486; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2488 = 10'h1b6 == ReadPtr[9:0] ? FifoCell_438 : _GEN_2487; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2489 = 10'h1b7 == ReadPtr[9:0] ? FifoCell_439 : _GEN_2488; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2490 = 10'h1b8 == ReadPtr[9:0] ? FifoCell_440 : _GEN_2489; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2491 = 10'h1b9 == ReadPtr[9:0] ? FifoCell_441 : _GEN_2490; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2492 = 10'h1ba == ReadPtr[9:0] ? FifoCell_442 : _GEN_2491; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2493 = 10'h1bb == ReadPtr[9:0] ? FifoCell_443 : _GEN_2492; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2494 = 10'h1bc == ReadPtr[9:0] ? FifoCell_444 : _GEN_2493; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2495 = 10'h1bd == ReadPtr[9:0] ? FifoCell_445 : _GEN_2494; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2496 = 10'h1be == ReadPtr[9:0] ? FifoCell_446 : _GEN_2495; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2497 = 10'h1bf == ReadPtr[9:0] ? FifoCell_447 : _GEN_2496; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2498 = 10'h1c0 == ReadPtr[9:0] ? FifoCell_448 : _GEN_2497; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2499 = 10'h1c1 == ReadPtr[9:0] ? FifoCell_449 : _GEN_2498; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2500 = 10'h1c2 == ReadPtr[9:0] ? FifoCell_450 : _GEN_2499; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2501 = 10'h1c3 == ReadPtr[9:0] ? FifoCell_451 : _GEN_2500; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2502 = 10'h1c4 == ReadPtr[9:0] ? FifoCell_452 : _GEN_2501; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2503 = 10'h1c5 == ReadPtr[9:0] ? FifoCell_453 : _GEN_2502; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2504 = 10'h1c6 == ReadPtr[9:0] ? FifoCell_454 : _GEN_2503; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2505 = 10'h1c7 == ReadPtr[9:0] ? FifoCell_455 : _GEN_2504; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2506 = 10'h1c8 == ReadPtr[9:0] ? FifoCell_456 : _GEN_2505; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2507 = 10'h1c9 == ReadPtr[9:0] ? FifoCell_457 : _GEN_2506; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2508 = 10'h1ca == ReadPtr[9:0] ? FifoCell_458 : _GEN_2507; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2509 = 10'h1cb == ReadPtr[9:0] ? FifoCell_459 : _GEN_2508; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2510 = 10'h1cc == ReadPtr[9:0] ? FifoCell_460 : _GEN_2509; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2511 = 10'h1cd == ReadPtr[9:0] ? FifoCell_461 : _GEN_2510; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2512 = 10'h1ce == ReadPtr[9:0] ? FifoCell_462 : _GEN_2511; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2513 = 10'h1cf == ReadPtr[9:0] ? FifoCell_463 : _GEN_2512; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2514 = 10'h1d0 == ReadPtr[9:0] ? FifoCell_464 : _GEN_2513; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2515 = 10'h1d1 == ReadPtr[9:0] ? FifoCell_465 : _GEN_2514; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2516 = 10'h1d2 == ReadPtr[9:0] ? FifoCell_466 : _GEN_2515; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2517 = 10'h1d3 == ReadPtr[9:0] ? FifoCell_467 : _GEN_2516; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2518 = 10'h1d4 == ReadPtr[9:0] ? FifoCell_468 : _GEN_2517; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2519 = 10'h1d5 == ReadPtr[9:0] ? FifoCell_469 : _GEN_2518; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2520 = 10'h1d6 == ReadPtr[9:0] ? FifoCell_470 : _GEN_2519; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2521 = 10'h1d7 == ReadPtr[9:0] ? FifoCell_471 : _GEN_2520; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2522 = 10'h1d8 == ReadPtr[9:0] ? FifoCell_472 : _GEN_2521; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2523 = 10'h1d9 == ReadPtr[9:0] ? FifoCell_473 : _GEN_2522; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2524 = 10'h1da == ReadPtr[9:0] ? FifoCell_474 : _GEN_2523; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2525 = 10'h1db == ReadPtr[9:0] ? FifoCell_475 : _GEN_2524; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2526 = 10'h1dc == ReadPtr[9:0] ? FifoCell_476 : _GEN_2525; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2527 = 10'h1dd == ReadPtr[9:0] ? FifoCell_477 : _GEN_2526; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2528 = 10'h1de == ReadPtr[9:0] ? FifoCell_478 : _GEN_2527; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2529 = 10'h1df == ReadPtr[9:0] ? FifoCell_479 : _GEN_2528; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2530 = 10'h1e0 == ReadPtr[9:0] ? FifoCell_480 : _GEN_2529; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2531 = 10'h1e1 == ReadPtr[9:0] ? FifoCell_481 : _GEN_2530; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2532 = 10'h1e2 == ReadPtr[9:0] ? FifoCell_482 : _GEN_2531; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2533 = 10'h1e3 == ReadPtr[9:0] ? FifoCell_483 : _GEN_2532; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2534 = 10'h1e4 == ReadPtr[9:0] ? FifoCell_484 : _GEN_2533; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2535 = 10'h1e5 == ReadPtr[9:0] ? FifoCell_485 : _GEN_2534; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2536 = 10'h1e6 == ReadPtr[9:0] ? FifoCell_486 : _GEN_2535; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2537 = 10'h1e7 == ReadPtr[9:0] ? FifoCell_487 : _GEN_2536; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2538 = 10'h1e8 == ReadPtr[9:0] ? FifoCell_488 : _GEN_2537; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2539 = 10'h1e9 == ReadPtr[9:0] ? FifoCell_489 : _GEN_2538; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2540 = 10'h1ea == ReadPtr[9:0] ? FifoCell_490 : _GEN_2539; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2541 = 10'h1eb == ReadPtr[9:0] ? FifoCell_491 : _GEN_2540; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2542 = 10'h1ec == ReadPtr[9:0] ? FifoCell_492 : _GEN_2541; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2543 = 10'h1ed == ReadPtr[9:0] ? FifoCell_493 : _GEN_2542; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2544 = 10'h1ee == ReadPtr[9:0] ? FifoCell_494 : _GEN_2543; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2545 = 10'h1ef == ReadPtr[9:0] ? FifoCell_495 : _GEN_2544; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2546 = 10'h1f0 == ReadPtr[9:0] ? FifoCell_496 : _GEN_2545; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2547 = 10'h1f1 == ReadPtr[9:0] ? FifoCell_497 : _GEN_2546; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2548 = 10'h1f2 == ReadPtr[9:0] ? FifoCell_498 : _GEN_2547; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2549 = 10'h1f3 == ReadPtr[9:0] ? FifoCell_499 : _GEN_2548; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2550 = 10'h1f4 == ReadPtr[9:0] ? FifoCell_500 : _GEN_2549; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2551 = 10'h1f5 == ReadPtr[9:0] ? FifoCell_501 : _GEN_2550; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2552 = 10'h1f6 == ReadPtr[9:0] ? FifoCell_502 : _GEN_2551; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2553 = 10'h1f7 == ReadPtr[9:0] ? FifoCell_503 : _GEN_2552; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2554 = 10'h1f8 == ReadPtr[9:0] ? FifoCell_504 : _GEN_2553; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2555 = 10'h1f9 == ReadPtr[9:0] ? FifoCell_505 : _GEN_2554; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2556 = 10'h1fa == ReadPtr[9:0] ? FifoCell_506 : _GEN_2555; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2557 = 10'h1fb == ReadPtr[9:0] ? FifoCell_507 : _GEN_2556; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2558 = 10'h1fc == ReadPtr[9:0] ? FifoCell_508 : _GEN_2557; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2559 = 10'h1fd == ReadPtr[9:0] ? FifoCell_509 : _GEN_2558; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2560 = 10'h1fe == ReadPtr[9:0] ? FifoCell_510 : _GEN_2559; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2561 = 10'h1ff == ReadPtr[9:0] ? FifoCell_511 : _GEN_2560; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2562 = 10'h200 == ReadPtr[9:0] ? FifoCell_512 : _GEN_2561; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2563 = 10'h201 == ReadPtr[9:0] ? FifoCell_513 : _GEN_2562; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2564 = 10'h202 == ReadPtr[9:0] ? FifoCell_514 : _GEN_2563; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2565 = 10'h203 == ReadPtr[9:0] ? FifoCell_515 : _GEN_2564; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2566 = 10'h204 == ReadPtr[9:0] ? FifoCell_516 : _GEN_2565; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2567 = 10'h205 == ReadPtr[9:0] ? FifoCell_517 : _GEN_2566; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2568 = 10'h206 == ReadPtr[9:0] ? FifoCell_518 : _GEN_2567; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2569 = 10'h207 == ReadPtr[9:0] ? FifoCell_519 : _GEN_2568; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2570 = 10'h208 == ReadPtr[9:0] ? FifoCell_520 : _GEN_2569; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2571 = 10'h209 == ReadPtr[9:0] ? FifoCell_521 : _GEN_2570; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2572 = 10'h20a == ReadPtr[9:0] ? FifoCell_522 : _GEN_2571; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2573 = 10'h20b == ReadPtr[9:0] ? FifoCell_523 : _GEN_2572; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2574 = 10'h20c == ReadPtr[9:0] ? FifoCell_524 : _GEN_2573; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2575 = 10'h20d == ReadPtr[9:0] ? FifoCell_525 : _GEN_2574; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2576 = 10'h20e == ReadPtr[9:0] ? FifoCell_526 : _GEN_2575; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2577 = 10'h20f == ReadPtr[9:0] ? FifoCell_527 : _GEN_2576; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2578 = 10'h210 == ReadPtr[9:0] ? FifoCell_528 : _GEN_2577; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2579 = 10'h211 == ReadPtr[9:0] ? FifoCell_529 : _GEN_2578; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2580 = 10'h212 == ReadPtr[9:0] ? FifoCell_530 : _GEN_2579; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2581 = 10'h213 == ReadPtr[9:0] ? FifoCell_531 : _GEN_2580; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2582 = 10'h214 == ReadPtr[9:0] ? FifoCell_532 : _GEN_2581; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2583 = 10'h215 == ReadPtr[9:0] ? FifoCell_533 : _GEN_2582; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2584 = 10'h216 == ReadPtr[9:0] ? FifoCell_534 : _GEN_2583; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2585 = 10'h217 == ReadPtr[9:0] ? FifoCell_535 : _GEN_2584; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2586 = 10'h218 == ReadPtr[9:0] ? FifoCell_536 : _GEN_2585; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2587 = 10'h219 == ReadPtr[9:0] ? FifoCell_537 : _GEN_2586; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2588 = 10'h21a == ReadPtr[9:0] ? FifoCell_538 : _GEN_2587; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2589 = 10'h21b == ReadPtr[9:0] ? FifoCell_539 : _GEN_2588; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2590 = 10'h21c == ReadPtr[9:0] ? FifoCell_540 : _GEN_2589; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2591 = 10'h21d == ReadPtr[9:0] ? FifoCell_541 : _GEN_2590; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2592 = 10'h21e == ReadPtr[9:0] ? FifoCell_542 : _GEN_2591; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2593 = 10'h21f == ReadPtr[9:0] ? FifoCell_543 : _GEN_2592; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2594 = 10'h220 == ReadPtr[9:0] ? FifoCell_544 : _GEN_2593; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2595 = 10'h221 == ReadPtr[9:0] ? FifoCell_545 : _GEN_2594; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2596 = 10'h222 == ReadPtr[9:0] ? FifoCell_546 : _GEN_2595; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2597 = 10'h223 == ReadPtr[9:0] ? FifoCell_547 : _GEN_2596; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2598 = 10'h224 == ReadPtr[9:0] ? FifoCell_548 : _GEN_2597; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2599 = 10'h225 == ReadPtr[9:0] ? FifoCell_549 : _GEN_2598; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2600 = 10'h226 == ReadPtr[9:0] ? FifoCell_550 : _GEN_2599; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2601 = 10'h227 == ReadPtr[9:0] ? FifoCell_551 : _GEN_2600; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2602 = 10'h228 == ReadPtr[9:0] ? FifoCell_552 : _GEN_2601; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2603 = 10'h229 == ReadPtr[9:0] ? FifoCell_553 : _GEN_2602; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2604 = 10'h22a == ReadPtr[9:0] ? FifoCell_554 : _GEN_2603; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2605 = 10'h22b == ReadPtr[9:0] ? FifoCell_555 : _GEN_2604; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2606 = 10'h22c == ReadPtr[9:0] ? FifoCell_556 : _GEN_2605; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2607 = 10'h22d == ReadPtr[9:0] ? FifoCell_557 : _GEN_2606; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2608 = 10'h22e == ReadPtr[9:0] ? FifoCell_558 : _GEN_2607; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2609 = 10'h22f == ReadPtr[9:0] ? FifoCell_559 : _GEN_2608; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2610 = 10'h230 == ReadPtr[9:0] ? FifoCell_560 : _GEN_2609; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2611 = 10'h231 == ReadPtr[9:0] ? FifoCell_561 : _GEN_2610; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2612 = 10'h232 == ReadPtr[9:0] ? FifoCell_562 : _GEN_2611; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2613 = 10'h233 == ReadPtr[9:0] ? FifoCell_563 : _GEN_2612; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2614 = 10'h234 == ReadPtr[9:0] ? FifoCell_564 : _GEN_2613; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2615 = 10'h235 == ReadPtr[9:0] ? FifoCell_565 : _GEN_2614; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2616 = 10'h236 == ReadPtr[9:0] ? FifoCell_566 : _GEN_2615; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2617 = 10'h237 == ReadPtr[9:0] ? FifoCell_567 : _GEN_2616; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2618 = 10'h238 == ReadPtr[9:0] ? FifoCell_568 : _GEN_2617; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2619 = 10'h239 == ReadPtr[9:0] ? FifoCell_569 : _GEN_2618; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2620 = 10'h23a == ReadPtr[9:0] ? FifoCell_570 : _GEN_2619; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2621 = 10'h23b == ReadPtr[9:0] ? FifoCell_571 : _GEN_2620; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2622 = 10'h23c == ReadPtr[9:0] ? FifoCell_572 : _GEN_2621; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2623 = 10'h23d == ReadPtr[9:0] ? FifoCell_573 : _GEN_2622; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2624 = 10'h23e == ReadPtr[9:0] ? FifoCell_574 : _GEN_2623; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2625 = 10'h23f == ReadPtr[9:0] ? FifoCell_575 : _GEN_2624; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2626 = 10'h240 == ReadPtr[9:0] ? FifoCell_576 : _GEN_2625; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2627 = 10'h241 == ReadPtr[9:0] ? FifoCell_577 : _GEN_2626; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2628 = 10'h242 == ReadPtr[9:0] ? FifoCell_578 : _GEN_2627; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2629 = 10'h243 == ReadPtr[9:0] ? FifoCell_579 : _GEN_2628; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2630 = 10'h244 == ReadPtr[9:0] ? FifoCell_580 : _GEN_2629; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2631 = 10'h245 == ReadPtr[9:0] ? FifoCell_581 : _GEN_2630; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2632 = 10'h246 == ReadPtr[9:0] ? FifoCell_582 : _GEN_2631; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2633 = 10'h247 == ReadPtr[9:0] ? FifoCell_583 : _GEN_2632; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2634 = 10'h248 == ReadPtr[9:0] ? FifoCell_584 : _GEN_2633; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2635 = 10'h249 == ReadPtr[9:0] ? FifoCell_585 : _GEN_2634; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2636 = 10'h24a == ReadPtr[9:0] ? FifoCell_586 : _GEN_2635; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2637 = 10'h24b == ReadPtr[9:0] ? FifoCell_587 : _GEN_2636; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2638 = 10'h24c == ReadPtr[9:0] ? FifoCell_588 : _GEN_2637; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2639 = 10'h24d == ReadPtr[9:0] ? FifoCell_589 : _GEN_2638; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2640 = 10'h24e == ReadPtr[9:0] ? FifoCell_590 : _GEN_2639; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2641 = 10'h24f == ReadPtr[9:0] ? FifoCell_591 : _GEN_2640; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2642 = 10'h250 == ReadPtr[9:0] ? FifoCell_592 : _GEN_2641; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2643 = 10'h251 == ReadPtr[9:0] ? FifoCell_593 : _GEN_2642; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2644 = 10'h252 == ReadPtr[9:0] ? FifoCell_594 : _GEN_2643; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2645 = 10'h253 == ReadPtr[9:0] ? FifoCell_595 : _GEN_2644; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2646 = 10'h254 == ReadPtr[9:0] ? FifoCell_596 : _GEN_2645; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2647 = 10'h255 == ReadPtr[9:0] ? FifoCell_597 : _GEN_2646; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2648 = 10'h256 == ReadPtr[9:0] ? FifoCell_598 : _GEN_2647; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2649 = 10'h257 == ReadPtr[9:0] ? FifoCell_599 : _GEN_2648; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2650 = 10'h258 == ReadPtr[9:0] ? FifoCell_600 : _GEN_2649; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2651 = 10'h259 == ReadPtr[9:0] ? FifoCell_601 : _GEN_2650; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2652 = 10'h25a == ReadPtr[9:0] ? FifoCell_602 : _GEN_2651; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2653 = 10'h25b == ReadPtr[9:0] ? FifoCell_603 : _GEN_2652; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2654 = 10'h25c == ReadPtr[9:0] ? FifoCell_604 : _GEN_2653; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2655 = 10'h25d == ReadPtr[9:0] ? FifoCell_605 : _GEN_2654; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2656 = 10'h25e == ReadPtr[9:0] ? FifoCell_606 : _GEN_2655; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2657 = 10'h25f == ReadPtr[9:0] ? FifoCell_607 : _GEN_2656; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2658 = 10'h260 == ReadPtr[9:0] ? FifoCell_608 : _GEN_2657; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2659 = 10'h261 == ReadPtr[9:0] ? FifoCell_609 : _GEN_2658; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2660 = 10'h262 == ReadPtr[9:0] ? FifoCell_610 : _GEN_2659; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2661 = 10'h263 == ReadPtr[9:0] ? FifoCell_611 : _GEN_2660; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2662 = 10'h264 == ReadPtr[9:0] ? FifoCell_612 : _GEN_2661; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2663 = 10'h265 == ReadPtr[9:0] ? FifoCell_613 : _GEN_2662; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2664 = 10'h266 == ReadPtr[9:0] ? FifoCell_614 : _GEN_2663; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2665 = 10'h267 == ReadPtr[9:0] ? FifoCell_615 : _GEN_2664; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2666 = 10'h268 == ReadPtr[9:0] ? FifoCell_616 : _GEN_2665; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2667 = 10'h269 == ReadPtr[9:0] ? FifoCell_617 : _GEN_2666; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2668 = 10'h26a == ReadPtr[9:0] ? FifoCell_618 : _GEN_2667; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2669 = 10'h26b == ReadPtr[9:0] ? FifoCell_619 : _GEN_2668; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2670 = 10'h26c == ReadPtr[9:0] ? FifoCell_620 : _GEN_2669; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2671 = 10'h26d == ReadPtr[9:0] ? FifoCell_621 : _GEN_2670; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2672 = 10'h26e == ReadPtr[9:0] ? FifoCell_622 : _GEN_2671; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2673 = 10'h26f == ReadPtr[9:0] ? FifoCell_623 : _GEN_2672; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2674 = 10'h270 == ReadPtr[9:0] ? FifoCell_624 : _GEN_2673; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2675 = 10'h271 == ReadPtr[9:0] ? FifoCell_625 : _GEN_2674; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2676 = 10'h272 == ReadPtr[9:0] ? FifoCell_626 : _GEN_2675; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2677 = 10'h273 == ReadPtr[9:0] ? FifoCell_627 : _GEN_2676; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2678 = 10'h274 == ReadPtr[9:0] ? FifoCell_628 : _GEN_2677; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2679 = 10'h275 == ReadPtr[9:0] ? FifoCell_629 : _GEN_2678; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2680 = 10'h276 == ReadPtr[9:0] ? FifoCell_630 : _GEN_2679; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2681 = 10'h277 == ReadPtr[9:0] ? FifoCell_631 : _GEN_2680; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2682 = 10'h278 == ReadPtr[9:0] ? FifoCell_632 : _GEN_2681; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2683 = 10'h279 == ReadPtr[9:0] ? FifoCell_633 : _GEN_2682; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2684 = 10'h27a == ReadPtr[9:0] ? FifoCell_634 : _GEN_2683; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2685 = 10'h27b == ReadPtr[9:0] ? FifoCell_635 : _GEN_2684; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2686 = 10'h27c == ReadPtr[9:0] ? FifoCell_636 : _GEN_2685; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2687 = 10'h27d == ReadPtr[9:0] ? FifoCell_637 : _GEN_2686; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2688 = 10'h27e == ReadPtr[9:0] ? FifoCell_638 : _GEN_2687; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2689 = 10'h27f == ReadPtr[9:0] ? FifoCell_639 : _GEN_2688; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2690 = 10'h280 == ReadPtr[9:0] ? FifoCell_640 : _GEN_2689; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2691 = 10'h281 == ReadPtr[9:0] ? FifoCell_641 : _GEN_2690; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2692 = 10'h282 == ReadPtr[9:0] ? FifoCell_642 : _GEN_2691; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2693 = 10'h283 == ReadPtr[9:0] ? FifoCell_643 : _GEN_2692; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2694 = 10'h284 == ReadPtr[9:0] ? FifoCell_644 : _GEN_2693; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2695 = 10'h285 == ReadPtr[9:0] ? FifoCell_645 : _GEN_2694; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2696 = 10'h286 == ReadPtr[9:0] ? FifoCell_646 : _GEN_2695; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2697 = 10'h287 == ReadPtr[9:0] ? FifoCell_647 : _GEN_2696; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2698 = 10'h288 == ReadPtr[9:0] ? FifoCell_648 : _GEN_2697; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2699 = 10'h289 == ReadPtr[9:0] ? FifoCell_649 : _GEN_2698; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2700 = 10'h28a == ReadPtr[9:0] ? FifoCell_650 : _GEN_2699; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2701 = 10'h28b == ReadPtr[9:0] ? FifoCell_651 : _GEN_2700; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2702 = 10'h28c == ReadPtr[9:0] ? FifoCell_652 : _GEN_2701; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2703 = 10'h28d == ReadPtr[9:0] ? FifoCell_653 : _GEN_2702; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2704 = 10'h28e == ReadPtr[9:0] ? FifoCell_654 : _GEN_2703; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2705 = 10'h28f == ReadPtr[9:0] ? FifoCell_655 : _GEN_2704; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2706 = 10'h290 == ReadPtr[9:0] ? FifoCell_656 : _GEN_2705; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2707 = 10'h291 == ReadPtr[9:0] ? FifoCell_657 : _GEN_2706; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2708 = 10'h292 == ReadPtr[9:0] ? FifoCell_658 : _GEN_2707; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2709 = 10'h293 == ReadPtr[9:0] ? FifoCell_659 : _GEN_2708; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2710 = 10'h294 == ReadPtr[9:0] ? FifoCell_660 : _GEN_2709; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2711 = 10'h295 == ReadPtr[9:0] ? FifoCell_661 : _GEN_2710; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2712 = 10'h296 == ReadPtr[9:0] ? FifoCell_662 : _GEN_2711; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2713 = 10'h297 == ReadPtr[9:0] ? FifoCell_663 : _GEN_2712; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2714 = 10'h298 == ReadPtr[9:0] ? FifoCell_664 : _GEN_2713; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2715 = 10'h299 == ReadPtr[9:0] ? FifoCell_665 : _GEN_2714; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2716 = 10'h29a == ReadPtr[9:0] ? FifoCell_666 : _GEN_2715; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2717 = 10'h29b == ReadPtr[9:0] ? FifoCell_667 : _GEN_2716; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2718 = 10'h29c == ReadPtr[9:0] ? FifoCell_668 : _GEN_2717; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2719 = 10'h29d == ReadPtr[9:0] ? FifoCell_669 : _GEN_2718; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2720 = 10'h29e == ReadPtr[9:0] ? FifoCell_670 : _GEN_2719; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2721 = 10'h29f == ReadPtr[9:0] ? FifoCell_671 : _GEN_2720; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2722 = 10'h2a0 == ReadPtr[9:0] ? FifoCell_672 : _GEN_2721; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2723 = 10'h2a1 == ReadPtr[9:0] ? FifoCell_673 : _GEN_2722; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2724 = 10'h2a2 == ReadPtr[9:0] ? FifoCell_674 : _GEN_2723; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2725 = 10'h2a3 == ReadPtr[9:0] ? FifoCell_675 : _GEN_2724; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2726 = 10'h2a4 == ReadPtr[9:0] ? FifoCell_676 : _GEN_2725; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2727 = 10'h2a5 == ReadPtr[9:0] ? FifoCell_677 : _GEN_2726; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2728 = 10'h2a6 == ReadPtr[9:0] ? FifoCell_678 : _GEN_2727; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2729 = 10'h2a7 == ReadPtr[9:0] ? FifoCell_679 : _GEN_2728; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2730 = 10'h2a8 == ReadPtr[9:0] ? FifoCell_680 : _GEN_2729; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2731 = 10'h2a9 == ReadPtr[9:0] ? FifoCell_681 : _GEN_2730; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2732 = 10'h2aa == ReadPtr[9:0] ? FifoCell_682 : _GEN_2731; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2733 = 10'h2ab == ReadPtr[9:0] ? FifoCell_683 : _GEN_2732; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2734 = 10'h2ac == ReadPtr[9:0] ? FifoCell_684 : _GEN_2733; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2735 = 10'h2ad == ReadPtr[9:0] ? FifoCell_685 : _GEN_2734; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2736 = 10'h2ae == ReadPtr[9:0] ? FifoCell_686 : _GEN_2735; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2737 = 10'h2af == ReadPtr[9:0] ? FifoCell_687 : _GEN_2736; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2738 = 10'h2b0 == ReadPtr[9:0] ? FifoCell_688 : _GEN_2737; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2739 = 10'h2b1 == ReadPtr[9:0] ? FifoCell_689 : _GEN_2738; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2740 = 10'h2b2 == ReadPtr[9:0] ? FifoCell_690 : _GEN_2739; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2741 = 10'h2b3 == ReadPtr[9:0] ? FifoCell_691 : _GEN_2740; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2742 = 10'h2b4 == ReadPtr[9:0] ? FifoCell_692 : _GEN_2741; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2743 = 10'h2b5 == ReadPtr[9:0] ? FifoCell_693 : _GEN_2742; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2744 = 10'h2b6 == ReadPtr[9:0] ? FifoCell_694 : _GEN_2743; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2745 = 10'h2b7 == ReadPtr[9:0] ? FifoCell_695 : _GEN_2744; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2746 = 10'h2b8 == ReadPtr[9:0] ? FifoCell_696 : _GEN_2745; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2747 = 10'h2b9 == ReadPtr[9:0] ? FifoCell_697 : _GEN_2746; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2748 = 10'h2ba == ReadPtr[9:0] ? FifoCell_698 : _GEN_2747; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2749 = 10'h2bb == ReadPtr[9:0] ? FifoCell_699 : _GEN_2748; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2750 = 10'h2bc == ReadPtr[9:0] ? FifoCell_700 : _GEN_2749; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2751 = 10'h2bd == ReadPtr[9:0] ? FifoCell_701 : _GEN_2750; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2752 = 10'h2be == ReadPtr[9:0] ? FifoCell_702 : _GEN_2751; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2753 = 10'h2bf == ReadPtr[9:0] ? FifoCell_703 : _GEN_2752; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2754 = 10'h2c0 == ReadPtr[9:0] ? FifoCell_704 : _GEN_2753; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2755 = 10'h2c1 == ReadPtr[9:0] ? FifoCell_705 : _GEN_2754; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2756 = 10'h2c2 == ReadPtr[9:0] ? FifoCell_706 : _GEN_2755; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2757 = 10'h2c3 == ReadPtr[9:0] ? FifoCell_707 : _GEN_2756; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2758 = 10'h2c4 == ReadPtr[9:0] ? FifoCell_708 : _GEN_2757; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2759 = 10'h2c5 == ReadPtr[9:0] ? FifoCell_709 : _GEN_2758; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2760 = 10'h2c6 == ReadPtr[9:0] ? FifoCell_710 : _GEN_2759; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2761 = 10'h2c7 == ReadPtr[9:0] ? FifoCell_711 : _GEN_2760; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2762 = 10'h2c8 == ReadPtr[9:0] ? FifoCell_712 : _GEN_2761; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2763 = 10'h2c9 == ReadPtr[9:0] ? FifoCell_713 : _GEN_2762; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2764 = 10'h2ca == ReadPtr[9:0] ? FifoCell_714 : _GEN_2763; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2765 = 10'h2cb == ReadPtr[9:0] ? FifoCell_715 : _GEN_2764; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2766 = 10'h2cc == ReadPtr[9:0] ? FifoCell_716 : _GEN_2765; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2767 = 10'h2cd == ReadPtr[9:0] ? FifoCell_717 : _GEN_2766; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2768 = 10'h2ce == ReadPtr[9:0] ? FifoCell_718 : _GEN_2767; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2769 = 10'h2cf == ReadPtr[9:0] ? FifoCell_719 : _GEN_2768; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2770 = 10'h2d0 == ReadPtr[9:0] ? FifoCell_720 : _GEN_2769; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2771 = 10'h2d1 == ReadPtr[9:0] ? FifoCell_721 : _GEN_2770; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2772 = 10'h2d2 == ReadPtr[9:0] ? FifoCell_722 : _GEN_2771; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2773 = 10'h2d3 == ReadPtr[9:0] ? FifoCell_723 : _GEN_2772; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2774 = 10'h2d4 == ReadPtr[9:0] ? FifoCell_724 : _GEN_2773; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2775 = 10'h2d5 == ReadPtr[9:0] ? FifoCell_725 : _GEN_2774; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2776 = 10'h2d6 == ReadPtr[9:0] ? FifoCell_726 : _GEN_2775; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2777 = 10'h2d7 == ReadPtr[9:0] ? FifoCell_727 : _GEN_2776; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2778 = 10'h2d8 == ReadPtr[9:0] ? FifoCell_728 : _GEN_2777; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2779 = 10'h2d9 == ReadPtr[9:0] ? FifoCell_729 : _GEN_2778; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2780 = 10'h2da == ReadPtr[9:0] ? FifoCell_730 : _GEN_2779; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2781 = 10'h2db == ReadPtr[9:0] ? FifoCell_731 : _GEN_2780; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2782 = 10'h2dc == ReadPtr[9:0] ? FifoCell_732 : _GEN_2781; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2783 = 10'h2dd == ReadPtr[9:0] ? FifoCell_733 : _GEN_2782; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2784 = 10'h2de == ReadPtr[9:0] ? FifoCell_734 : _GEN_2783; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2785 = 10'h2df == ReadPtr[9:0] ? FifoCell_735 : _GEN_2784; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2786 = 10'h2e0 == ReadPtr[9:0] ? FifoCell_736 : _GEN_2785; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2787 = 10'h2e1 == ReadPtr[9:0] ? FifoCell_737 : _GEN_2786; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2788 = 10'h2e2 == ReadPtr[9:0] ? FifoCell_738 : _GEN_2787; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2789 = 10'h2e3 == ReadPtr[9:0] ? FifoCell_739 : _GEN_2788; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2790 = 10'h2e4 == ReadPtr[9:0] ? FifoCell_740 : _GEN_2789; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2791 = 10'h2e5 == ReadPtr[9:0] ? FifoCell_741 : _GEN_2790; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2792 = 10'h2e6 == ReadPtr[9:0] ? FifoCell_742 : _GEN_2791; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2793 = 10'h2e7 == ReadPtr[9:0] ? FifoCell_743 : _GEN_2792; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2794 = 10'h2e8 == ReadPtr[9:0] ? FifoCell_744 : _GEN_2793; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2795 = 10'h2e9 == ReadPtr[9:0] ? FifoCell_745 : _GEN_2794; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2796 = 10'h2ea == ReadPtr[9:0] ? FifoCell_746 : _GEN_2795; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2797 = 10'h2eb == ReadPtr[9:0] ? FifoCell_747 : _GEN_2796; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2798 = 10'h2ec == ReadPtr[9:0] ? FifoCell_748 : _GEN_2797; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2799 = 10'h2ed == ReadPtr[9:0] ? FifoCell_749 : _GEN_2798; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2800 = 10'h2ee == ReadPtr[9:0] ? FifoCell_750 : _GEN_2799; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2801 = 10'h2ef == ReadPtr[9:0] ? FifoCell_751 : _GEN_2800; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2802 = 10'h2f0 == ReadPtr[9:0] ? FifoCell_752 : _GEN_2801; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2803 = 10'h2f1 == ReadPtr[9:0] ? FifoCell_753 : _GEN_2802; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2804 = 10'h2f2 == ReadPtr[9:0] ? FifoCell_754 : _GEN_2803; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2805 = 10'h2f3 == ReadPtr[9:0] ? FifoCell_755 : _GEN_2804; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2806 = 10'h2f4 == ReadPtr[9:0] ? FifoCell_756 : _GEN_2805; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2807 = 10'h2f5 == ReadPtr[9:0] ? FifoCell_757 : _GEN_2806; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2808 = 10'h2f6 == ReadPtr[9:0] ? FifoCell_758 : _GEN_2807; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2809 = 10'h2f7 == ReadPtr[9:0] ? FifoCell_759 : _GEN_2808; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2810 = 10'h2f8 == ReadPtr[9:0] ? FifoCell_760 : _GEN_2809; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2811 = 10'h2f9 == ReadPtr[9:0] ? FifoCell_761 : _GEN_2810; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2812 = 10'h2fa == ReadPtr[9:0] ? FifoCell_762 : _GEN_2811; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2813 = 10'h2fb == ReadPtr[9:0] ? FifoCell_763 : _GEN_2812; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2814 = 10'h2fc == ReadPtr[9:0] ? FifoCell_764 : _GEN_2813; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2815 = 10'h2fd == ReadPtr[9:0] ? FifoCell_765 : _GEN_2814; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2816 = 10'h2fe == ReadPtr[9:0] ? FifoCell_766 : _GEN_2815; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2817 = 10'h2ff == ReadPtr[9:0] ? FifoCell_767 : _GEN_2816; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2818 = 10'h300 == ReadPtr[9:0] ? FifoCell_768 : _GEN_2817; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2819 = 10'h301 == ReadPtr[9:0] ? FifoCell_769 : _GEN_2818; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2820 = 10'h302 == ReadPtr[9:0] ? FifoCell_770 : _GEN_2819; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2821 = 10'h303 == ReadPtr[9:0] ? FifoCell_771 : _GEN_2820; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2822 = 10'h304 == ReadPtr[9:0] ? FifoCell_772 : _GEN_2821; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2823 = 10'h305 == ReadPtr[9:0] ? FifoCell_773 : _GEN_2822; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2824 = 10'h306 == ReadPtr[9:0] ? FifoCell_774 : _GEN_2823; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2825 = 10'h307 == ReadPtr[9:0] ? FifoCell_775 : _GEN_2824; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2826 = 10'h308 == ReadPtr[9:0] ? FifoCell_776 : _GEN_2825; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2827 = 10'h309 == ReadPtr[9:0] ? FifoCell_777 : _GEN_2826; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2828 = 10'h30a == ReadPtr[9:0] ? FifoCell_778 : _GEN_2827; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2829 = 10'h30b == ReadPtr[9:0] ? FifoCell_779 : _GEN_2828; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2830 = 10'h30c == ReadPtr[9:0] ? FifoCell_780 : _GEN_2829; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2831 = 10'h30d == ReadPtr[9:0] ? FifoCell_781 : _GEN_2830; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2832 = 10'h30e == ReadPtr[9:0] ? FifoCell_782 : _GEN_2831; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2833 = 10'h30f == ReadPtr[9:0] ? FifoCell_783 : _GEN_2832; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2834 = 10'h310 == ReadPtr[9:0] ? FifoCell_784 : _GEN_2833; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2835 = 10'h311 == ReadPtr[9:0] ? FifoCell_785 : _GEN_2834; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2836 = 10'h312 == ReadPtr[9:0] ? FifoCell_786 : _GEN_2835; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2837 = 10'h313 == ReadPtr[9:0] ? FifoCell_787 : _GEN_2836; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2838 = 10'h314 == ReadPtr[9:0] ? FifoCell_788 : _GEN_2837; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2839 = 10'h315 == ReadPtr[9:0] ? FifoCell_789 : _GEN_2838; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2840 = 10'h316 == ReadPtr[9:0] ? FifoCell_790 : _GEN_2839; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2841 = 10'h317 == ReadPtr[9:0] ? FifoCell_791 : _GEN_2840; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2842 = 10'h318 == ReadPtr[9:0] ? FifoCell_792 : _GEN_2841; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2843 = 10'h319 == ReadPtr[9:0] ? FifoCell_793 : _GEN_2842; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2844 = 10'h31a == ReadPtr[9:0] ? FifoCell_794 : _GEN_2843; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2845 = 10'h31b == ReadPtr[9:0] ? FifoCell_795 : _GEN_2844; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2846 = 10'h31c == ReadPtr[9:0] ? FifoCell_796 : _GEN_2845; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2847 = 10'h31d == ReadPtr[9:0] ? FifoCell_797 : _GEN_2846; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2848 = 10'h31e == ReadPtr[9:0] ? FifoCell_798 : _GEN_2847; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2849 = 10'h31f == ReadPtr[9:0] ? FifoCell_799 : _GEN_2848; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2850 = 10'h320 == ReadPtr[9:0] ? FifoCell_800 : _GEN_2849; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2851 = 10'h321 == ReadPtr[9:0] ? FifoCell_801 : _GEN_2850; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2852 = 10'h322 == ReadPtr[9:0] ? FifoCell_802 : _GEN_2851; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2853 = 10'h323 == ReadPtr[9:0] ? FifoCell_803 : _GEN_2852; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2854 = 10'h324 == ReadPtr[9:0] ? FifoCell_804 : _GEN_2853; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2855 = 10'h325 == ReadPtr[9:0] ? FifoCell_805 : _GEN_2854; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2856 = 10'h326 == ReadPtr[9:0] ? FifoCell_806 : _GEN_2855; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2857 = 10'h327 == ReadPtr[9:0] ? FifoCell_807 : _GEN_2856; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2858 = 10'h328 == ReadPtr[9:0] ? FifoCell_808 : _GEN_2857; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2859 = 10'h329 == ReadPtr[9:0] ? FifoCell_809 : _GEN_2858; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2860 = 10'h32a == ReadPtr[9:0] ? FifoCell_810 : _GEN_2859; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2861 = 10'h32b == ReadPtr[9:0] ? FifoCell_811 : _GEN_2860; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2862 = 10'h32c == ReadPtr[9:0] ? FifoCell_812 : _GEN_2861; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2863 = 10'h32d == ReadPtr[9:0] ? FifoCell_813 : _GEN_2862; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2864 = 10'h32e == ReadPtr[9:0] ? FifoCell_814 : _GEN_2863; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2865 = 10'h32f == ReadPtr[9:0] ? FifoCell_815 : _GEN_2864; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2866 = 10'h330 == ReadPtr[9:0] ? FifoCell_816 : _GEN_2865; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2867 = 10'h331 == ReadPtr[9:0] ? FifoCell_817 : _GEN_2866; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2868 = 10'h332 == ReadPtr[9:0] ? FifoCell_818 : _GEN_2867; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2869 = 10'h333 == ReadPtr[9:0] ? FifoCell_819 : _GEN_2868; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2870 = 10'h334 == ReadPtr[9:0] ? FifoCell_820 : _GEN_2869; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2871 = 10'h335 == ReadPtr[9:0] ? FifoCell_821 : _GEN_2870; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2872 = 10'h336 == ReadPtr[9:0] ? FifoCell_822 : _GEN_2871; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2873 = 10'h337 == ReadPtr[9:0] ? FifoCell_823 : _GEN_2872; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2874 = 10'h338 == ReadPtr[9:0] ? FifoCell_824 : _GEN_2873; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2875 = 10'h339 == ReadPtr[9:0] ? FifoCell_825 : _GEN_2874; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2876 = 10'h33a == ReadPtr[9:0] ? FifoCell_826 : _GEN_2875; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2877 = 10'h33b == ReadPtr[9:0] ? FifoCell_827 : _GEN_2876; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2878 = 10'h33c == ReadPtr[9:0] ? FifoCell_828 : _GEN_2877; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2879 = 10'h33d == ReadPtr[9:0] ? FifoCell_829 : _GEN_2878; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2880 = 10'h33e == ReadPtr[9:0] ? FifoCell_830 : _GEN_2879; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2881 = 10'h33f == ReadPtr[9:0] ? FifoCell_831 : _GEN_2880; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2882 = 10'h340 == ReadPtr[9:0] ? FifoCell_832 : _GEN_2881; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2883 = 10'h341 == ReadPtr[9:0] ? FifoCell_833 : _GEN_2882; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2884 = 10'h342 == ReadPtr[9:0] ? FifoCell_834 : _GEN_2883; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2885 = 10'h343 == ReadPtr[9:0] ? FifoCell_835 : _GEN_2884; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2886 = 10'h344 == ReadPtr[9:0] ? FifoCell_836 : _GEN_2885; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2887 = 10'h345 == ReadPtr[9:0] ? FifoCell_837 : _GEN_2886; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2888 = 10'h346 == ReadPtr[9:0] ? FifoCell_838 : _GEN_2887; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2889 = 10'h347 == ReadPtr[9:0] ? FifoCell_839 : _GEN_2888; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2890 = 10'h348 == ReadPtr[9:0] ? FifoCell_840 : _GEN_2889; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2891 = 10'h349 == ReadPtr[9:0] ? FifoCell_841 : _GEN_2890; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2892 = 10'h34a == ReadPtr[9:0] ? FifoCell_842 : _GEN_2891; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2893 = 10'h34b == ReadPtr[9:0] ? FifoCell_843 : _GEN_2892; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2894 = 10'h34c == ReadPtr[9:0] ? FifoCell_844 : _GEN_2893; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2895 = 10'h34d == ReadPtr[9:0] ? FifoCell_845 : _GEN_2894; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2896 = 10'h34e == ReadPtr[9:0] ? FifoCell_846 : _GEN_2895; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2897 = 10'h34f == ReadPtr[9:0] ? FifoCell_847 : _GEN_2896; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2898 = 10'h350 == ReadPtr[9:0] ? FifoCell_848 : _GEN_2897; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2899 = 10'h351 == ReadPtr[9:0] ? FifoCell_849 : _GEN_2898; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2900 = 10'h352 == ReadPtr[9:0] ? FifoCell_850 : _GEN_2899; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2901 = 10'h353 == ReadPtr[9:0] ? FifoCell_851 : _GEN_2900; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2902 = 10'h354 == ReadPtr[9:0] ? FifoCell_852 : _GEN_2901; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2903 = 10'h355 == ReadPtr[9:0] ? FifoCell_853 : _GEN_2902; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2904 = 10'h356 == ReadPtr[9:0] ? FifoCell_854 : _GEN_2903; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2905 = 10'h357 == ReadPtr[9:0] ? FifoCell_855 : _GEN_2904; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2906 = 10'h358 == ReadPtr[9:0] ? FifoCell_856 : _GEN_2905; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2907 = 10'h359 == ReadPtr[9:0] ? FifoCell_857 : _GEN_2906; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2908 = 10'h35a == ReadPtr[9:0] ? FifoCell_858 : _GEN_2907; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2909 = 10'h35b == ReadPtr[9:0] ? FifoCell_859 : _GEN_2908; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2910 = 10'h35c == ReadPtr[9:0] ? FifoCell_860 : _GEN_2909; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2911 = 10'h35d == ReadPtr[9:0] ? FifoCell_861 : _GEN_2910; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2912 = 10'h35e == ReadPtr[9:0] ? FifoCell_862 : _GEN_2911; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2913 = 10'h35f == ReadPtr[9:0] ? FifoCell_863 : _GEN_2912; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2914 = 10'h360 == ReadPtr[9:0] ? FifoCell_864 : _GEN_2913; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2915 = 10'h361 == ReadPtr[9:0] ? FifoCell_865 : _GEN_2914; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2916 = 10'h362 == ReadPtr[9:0] ? FifoCell_866 : _GEN_2915; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2917 = 10'h363 == ReadPtr[9:0] ? FifoCell_867 : _GEN_2916; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2918 = 10'h364 == ReadPtr[9:0] ? FifoCell_868 : _GEN_2917; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2919 = 10'h365 == ReadPtr[9:0] ? FifoCell_869 : _GEN_2918; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2920 = 10'h366 == ReadPtr[9:0] ? FifoCell_870 : _GEN_2919; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2921 = 10'h367 == ReadPtr[9:0] ? FifoCell_871 : _GEN_2920; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2922 = 10'h368 == ReadPtr[9:0] ? FifoCell_872 : _GEN_2921; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2923 = 10'h369 == ReadPtr[9:0] ? FifoCell_873 : _GEN_2922; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2924 = 10'h36a == ReadPtr[9:0] ? FifoCell_874 : _GEN_2923; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2925 = 10'h36b == ReadPtr[9:0] ? FifoCell_875 : _GEN_2924; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2926 = 10'h36c == ReadPtr[9:0] ? FifoCell_876 : _GEN_2925; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2927 = 10'h36d == ReadPtr[9:0] ? FifoCell_877 : _GEN_2926; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2928 = 10'h36e == ReadPtr[9:0] ? FifoCell_878 : _GEN_2927; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2929 = 10'h36f == ReadPtr[9:0] ? FifoCell_879 : _GEN_2928; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2930 = 10'h370 == ReadPtr[9:0] ? FifoCell_880 : _GEN_2929; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2931 = 10'h371 == ReadPtr[9:0] ? FifoCell_881 : _GEN_2930; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2932 = 10'h372 == ReadPtr[9:0] ? FifoCell_882 : _GEN_2931; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2933 = 10'h373 == ReadPtr[9:0] ? FifoCell_883 : _GEN_2932; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2934 = 10'h374 == ReadPtr[9:0] ? FifoCell_884 : _GEN_2933; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2935 = 10'h375 == ReadPtr[9:0] ? FifoCell_885 : _GEN_2934; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2936 = 10'h376 == ReadPtr[9:0] ? FifoCell_886 : _GEN_2935; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2937 = 10'h377 == ReadPtr[9:0] ? FifoCell_887 : _GEN_2936; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2938 = 10'h378 == ReadPtr[9:0] ? FifoCell_888 : _GEN_2937; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2939 = 10'h379 == ReadPtr[9:0] ? FifoCell_889 : _GEN_2938; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2940 = 10'h37a == ReadPtr[9:0] ? FifoCell_890 : _GEN_2939; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2941 = 10'h37b == ReadPtr[9:0] ? FifoCell_891 : _GEN_2940; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2942 = 10'h37c == ReadPtr[9:0] ? FifoCell_892 : _GEN_2941; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2943 = 10'h37d == ReadPtr[9:0] ? FifoCell_893 : _GEN_2942; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2944 = 10'h37e == ReadPtr[9:0] ? FifoCell_894 : _GEN_2943; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2945 = 10'h37f == ReadPtr[9:0] ? FifoCell_895 : _GEN_2944; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2946 = 10'h380 == ReadPtr[9:0] ? FifoCell_896 : _GEN_2945; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2947 = 10'h381 == ReadPtr[9:0] ? FifoCell_897 : _GEN_2946; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2948 = 10'h382 == ReadPtr[9:0] ? FifoCell_898 : _GEN_2947; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2949 = 10'h383 == ReadPtr[9:0] ? FifoCell_899 : _GEN_2948; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2950 = 10'h384 == ReadPtr[9:0] ? FifoCell_900 : _GEN_2949; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2951 = 10'h385 == ReadPtr[9:0] ? FifoCell_901 : _GEN_2950; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2952 = 10'h386 == ReadPtr[9:0] ? FifoCell_902 : _GEN_2951; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2953 = 10'h387 == ReadPtr[9:0] ? FifoCell_903 : _GEN_2952; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2954 = 10'h388 == ReadPtr[9:0] ? FifoCell_904 : _GEN_2953; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2955 = 10'h389 == ReadPtr[9:0] ? FifoCell_905 : _GEN_2954; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2956 = 10'h38a == ReadPtr[9:0] ? FifoCell_906 : _GEN_2955; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2957 = 10'h38b == ReadPtr[9:0] ? FifoCell_907 : _GEN_2956; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2958 = 10'h38c == ReadPtr[9:0] ? FifoCell_908 : _GEN_2957; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2959 = 10'h38d == ReadPtr[9:0] ? FifoCell_909 : _GEN_2958; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2960 = 10'h38e == ReadPtr[9:0] ? FifoCell_910 : _GEN_2959; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2961 = 10'h38f == ReadPtr[9:0] ? FifoCell_911 : _GEN_2960; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2962 = 10'h390 == ReadPtr[9:0] ? FifoCell_912 : _GEN_2961; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2963 = 10'h391 == ReadPtr[9:0] ? FifoCell_913 : _GEN_2962; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2964 = 10'h392 == ReadPtr[9:0] ? FifoCell_914 : _GEN_2963; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2965 = 10'h393 == ReadPtr[9:0] ? FifoCell_915 : _GEN_2964; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2966 = 10'h394 == ReadPtr[9:0] ? FifoCell_916 : _GEN_2965; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2967 = 10'h395 == ReadPtr[9:0] ? FifoCell_917 : _GEN_2966; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2968 = 10'h396 == ReadPtr[9:0] ? FifoCell_918 : _GEN_2967; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2969 = 10'h397 == ReadPtr[9:0] ? FifoCell_919 : _GEN_2968; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2970 = 10'h398 == ReadPtr[9:0] ? FifoCell_920 : _GEN_2969; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2971 = 10'h399 == ReadPtr[9:0] ? FifoCell_921 : _GEN_2970; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2972 = 10'h39a == ReadPtr[9:0] ? FifoCell_922 : _GEN_2971; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2973 = 10'h39b == ReadPtr[9:0] ? FifoCell_923 : _GEN_2972; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2974 = 10'h39c == ReadPtr[9:0] ? FifoCell_924 : _GEN_2973; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2975 = 10'h39d == ReadPtr[9:0] ? FifoCell_925 : _GEN_2974; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2976 = 10'h39e == ReadPtr[9:0] ? FifoCell_926 : _GEN_2975; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2977 = 10'h39f == ReadPtr[9:0] ? FifoCell_927 : _GEN_2976; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2978 = 10'h3a0 == ReadPtr[9:0] ? FifoCell_928 : _GEN_2977; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2979 = 10'h3a1 == ReadPtr[9:0] ? FifoCell_929 : _GEN_2978; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2980 = 10'h3a2 == ReadPtr[9:0] ? FifoCell_930 : _GEN_2979; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2981 = 10'h3a3 == ReadPtr[9:0] ? FifoCell_931 : _GEN_2980; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2982 = 10'h3a4 == ReadPtr[9:0] ? FifoCell_932 : _GEN_2981; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2983 = 10'h3a5 == ReadPtr[9:0] ? FifoCell_933 : _GEN_2982; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2984 = 10'h3a6 == ReadPtr[9:0] ? FifoCell_934 : _GEN_2983; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2985 = 10'h3a7 == ReadPtr[9:0] ? FifoCell_935 : _GEN_2984; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2986 = 10'h3a8 == ReadPtr[9:0] ? FifoCell_936 : _GEN_2985; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2987 = 10'h3a9 == ReadPtr[9:0] ? FifoCell_937 : _GEN_2986; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2988 = 10'h3aa == ReadPtr[9:0] ? FifoCell_938 : _GEN_2987; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2989 = 10'h3ab == ReadPtr[9:0] ? FifoCell_939 : _GEN_2988; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2990 = 10'h3ac == ReadPtr[9:0] ? FifoCell_940 : _GEN_2989; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2991 = 10'h3ad == ReadPtr[9:0] ? FifoCell_941 : _GEN_2990; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2992 = 10'h3ae == ReadPtr[9:0] ? FifoCell_942 : _GEN_2991; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2993 = 10'h3af == ReadPtr[9:0] ? FifoCell_943 : _GEN_2992; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2994 = 10'h3b0 == ReadPtr[9:0] ? FifoCell_944 : _GEN_2993; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2995 = 10'h3b1 == ReadPtr[9:0] ? FifoCell_945 : _GEN_2994; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2996 = 10'h3b2 == ReadPtr[9:0] ? FifoCell_946 : _GEN_2995; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2997 = 10'h3b3 == ReadPtr[9:0] ? FifoCell_947 : _GEN_2996; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2998 = 10'h3b4 == ReadPtr[9:0] ? FifoCell_948 : _GEN_2997; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_2999 = 10'h3b5 == ReadPtr[9:0] ? FifoCell_949 : _GEN_2998; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_3000 = 10'h3b6 == ReadPtr[9:0] ? FifoCell_950 : _GEN_2999; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_3001 = 10'h3b7 == ReadPtr[9:0] ? FifoCell_951 : _GEN_3000; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_3002 = 10'h3b8 == ReadPtr[9:0] ? FifoCell_952 : _GEN_3001; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_3003 = 10'h3b9 == ReadPtr[9:0] ? FifoCell_953 : _GEN_3002; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_3004 = 10'h3ba == ReadPtr[9:0] ? FifoCell_954 : _GEN_3003; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_3005 = 10'h3bb == ReadPtr[9:0] ? FifoCell_955 : _GEN_3004; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_3006 = 10'h3bc == ReadPtr[9:0] ? FifoCell_956 : _GEN_3005; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_3007 = 10'h3bd == ReadPtr[9:0] ? FifoCell_957 : _GEN_3006; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_3008 = 10'h3be == ReadPtr[9:0] ? FifoCell_958 : _GEN_3007; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_3009 = 10'h3bf == ReadPtr[9:0] ? FifoCell_959 : _GEN_3008; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_3010 = 10'h3c0 == ReadPtr[9:0] ? FifoCell_960 : _GEN_3009; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_3011 = 10'h3c1 == ReadPtr[9:0] ? FifoCell_961 : _GEN_3010; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_3012 = 10'h3c2 == ReadPtr[9:0] ? FifoCell_962 : _GEN_3011; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_3013 = 10'h3c3 == ReadPtr[9:0] ? FifoCell_963 : _GEN_3012; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_3014 = 10'h3c4 == ReadPtr[9:0] ? FifoCell_964 : _GEN_3013; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_3015 = 10'h3c5 == ReadPtr[9:0] ? FifoCell_965 : _GEN_3014; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_3016 = 10'h3c6 == ReadPtr[9:0] ? FifoCell_966 : _GEN_3015; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_3017 = 10'h3c7 == ReadPtr[9:0] ? FifoCell_967 : _GEN_3016; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_3018 = 10'h3c8 == ReadPtr[9:0] ? FifoCell_968 : _GEN_3017; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_3019 = 10'h3c9 == ReadPtr[9:0] ? FifoCell_969 : _GEN_3018; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_3020 = 10'h3ca == ReadPtr[9:0] ? FifoCell_970 : _GEN_3019; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_3021 = 10'h3cb == ReadPtr[9:0] ? FifoCell_971 : _GEN_3020; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_3022 = 10'h3cc == ReadPtr[9:0] ? FifoCell_972 : _GEN_3021; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_3023 = 10'h3cd == ReadPtr[9:0] ? FifoCell_973 : _GEN_3022; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_3024 = 10'h3ce == ReadPtr[9:0] ? FifoCell_974 : _GEN_3023; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_3025 = 10'h3cf == ReadPtr[9:0] ? FifoCell_975 : _GEN_3024; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_3026 = 10'h3d0 == ReadPtr[9:0] ? FifoCell_976 : _GEN_3025; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_3027 = 10'h3d1 == ReadPtr[9:0] ? FifoCell_977 : _GEN_3026; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_3028 = 10'h3d2 == ReadPtr[9:0] ? FifoCell_978 : _GEN_3027; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_3029 = 10'h3d3 == ReadPtr[9:0] ? FifoCell_979 : _GEN_3028; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_3030 = 10'h3d4 == ReadPtr[9:0] ? FifoCell_980 : _GEN_3029; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_3031 = 10'h3d5 == ReadPtr[9:0] ? FifoCell_981 : _GEN_3030; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_3032 = 10'h3d6 == ReadPtr[9:0] ? FifoCell_982 : _GEN_3031; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_3033 = 10'h3d7 == ReadPtr[9:0] ? FifoCell_983 : _GEN_3032; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_3034 = 10'h3d8 == ReadPtr[9:0] ? FifoCell_984 : _GEN_3033; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_3035 = 10'h3d9 == ReadPtr[9:0] ? FifoCell_985 : _GEN_3034; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_3036 = 10'h3da == ReadPtr[9:0] ? FifoCell_986 : _GEN_3035; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_3037 = 10'h3db == ReadPtr[9:0] ? FifoCell_987 : _GEN_3036; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_3038 = 10'h3dc == ReadPtr[9:0] ? FifoCell_988 : _GEN_3037; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_3039 = 10'h3dd == ReadPtr[9:0] ? FifoCell_989 : _GEN_3038; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_3040 = 10'h3de == ReadPtr[9:0] ? FifoCell_990 : _GEN_3039; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_3041 = 10'h3df == ReadPtr[9:0] ? FifoCell_991 : _GEN_3040; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_3042 = 10'h3e0 == ReadPtr[9:0] ? FifoCell_992 : _GEN_3041; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_3043 = 10'h3e1 == ReadPtr[9:0] ? FifoCell_993 : _GEN_3042; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_3044 = 10'h3e2 == ReadPtr[9:0] ? FifoCell_994 : _GEN_3043; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_3045 = 10'h3e3 == ReadPtr[9:0] ? FifoCell_995 : _GEN_3044; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_3046 = 10'h3e4 == ReadPtr[9:0] ? FifoCell_996 : _GEN_3045; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_3047 = 10'h3e5 == ReadPtr[9:0] ? FifoCell_997 : _GEN_3046; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_3048 = 10'h3e6 == ReadPtr[9:0] ? FifoCell_998 : _GEN_3047; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_3049 = 10'h3e7 == ReadPtr[9:0] ? FifoCell_999 : _GEN_3048; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_3050 = 10'h3e8 == ReadPtr[9:0] ? FifoCell_1000 : _GEN_3049; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_3051 = 10'h3e9 == ReadPtr[9:0] ? FifoCell_1001 : _GEN_3050; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_3052 = 10'h3ea == ReadPtr[9:0] ? FifoCell_1002 : _GEN_3051; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_3053 = 10'h3eb == ReadPtr[9:0] ? FifoCell_1003 : _GEN_3052; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_3054 = 10'h3ec == ReadPtr[9:0] ? FifoCell_1004 : _GEN_3053; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_3055 = 10'h3ed == ReadPtr[9:0] ? FifoCell_1005 : _GEN_3054; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_3056 = 10'h3ee == ReadPtr[9:0] ? FifoCell_1006 : _GEN_3055; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_3057 = 10'h3ef == ReadPtr[9:0] ? FifoCell_1007 : _GEN_3056; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_3058 = 10'h3f0 == ReadPtr[9:0] ? FifoCell_1008 : _GEN_3057; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_3059 = 10'h3f1 == ReadPtr[9:0] ? FifoCell_1009 : _GEN_3058; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_3060 = 10'h3f2 == ReadPtr[9:0] ? FifoCell_1010 : _GEN_3059; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_3061 = 10'h3f3 == ReadPtr[9:0] ? FifoCell_1011 : _GEN_3060; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_3062 = 10'h3f4 == ReadPtr[9:0] ? FifoCell_1012 : _GEN_3061; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_3063 = 10'h3f5 == ReadPtr[9:0] ? FifoCell_1013 : _GEN_3062; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_3064 = 10'h3f6 == ReadPtr[9:0] ? FifoCell_1014 : _GEN_3063; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_3065 = 10'h3f7 == ReadPtr[9:0] ? FifoCell_1015 : _GEN_3064; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_3066 = 10'h3f8 == ReadPtr[9:0] ? FifoCell_1016 : _GEN_3065; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_3067 = 10'h3f9 == ReadPtr[9:0] ? FifoCell_1017 : _GEN_3066; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_3068 = 10'h3fa == ReadPtr[9:0] ? FifoCell_1018 : _GEN_3067; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_3069 = 10'h3fb == ReadPtr[9:0] ? FifoCell_1019 : _GEN_3068; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_3070 = 10'h3fc == ReadPtr[9:0] ? FifoCell_1020 : _GEN_3069; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_3071 = 10'h3fd == ReadPtr[9:0] ? FifoCell_1021 : _GEN_3070; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  wire [8:0] _GEN_3072 = 10'h3fe == ReadPtr[9:0] ? FifoCell_1022 : _GEN_3071; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  assign io_Writer_Full = WritePtr[10] != ReadPtr[10] & _io_Writer_Full_T_5; // @[src/main/scala/fifo_pkg/FifoPkg.scala 30:80]
  assign io_Reader_ReadData = 10'h3ff == ReadPtr[9:0] ? FifoCell_1023 : _GEN_3072; // @[src/main/scala/fifo_pkg/FifoPkg.scala 46:{22,22}]
  assign io_Reader_Empty = WritePtr == ReadPtr; // @[src/main/scala/fifo_pkg/FifoPkg.scala 32:32]
  always @(posedge clock) begin
    if (reset) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 26:25]
      WritePtr <= 11'h0; // @[src/main/scala/fifo_pkg/FifoPkg.scala 26:25]
    end else if (~io_Writer_Full & io_Writer_WriteEn) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 34:62]
      WritePtr <= _WritePtr_T_1; // @[src/main/scala/fifo_pkg/FifoPkg.scala 35:14]
    end
    if (reset) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 27:24]
      ReadPtr <= 11'h0; // @[src/main/scala/fifo_pkg/FifoPkg.scala 27:24]
    end else if (~io_Reader_Empty & io_Reader_ReadEn) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 38:62]
      ReadPtr <= _ReadPtr_T_1; // @[src/main/scala/fifo_pkg/FifoPkg.scala 39:13]
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h0 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_0 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h1 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_1 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h2 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_2 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h3 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_3 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h4 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_4 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h5 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_5 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h6 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_6 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h7 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_7 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h8 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_8 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h9 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_9 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'ha == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_10 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'hb == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_11 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'hc == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_12 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'hd == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_13 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'he == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_14 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'hf == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_15 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h10 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_16 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h11 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_17 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h12 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_18 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h13 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_19 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h14 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_20 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h15 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_21 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h16 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_22 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h17 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_23 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h18 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_24 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h19 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_25 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h1a == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_26 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h1b == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_27 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h1c == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_28 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h1d == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_29 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h1e == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_30 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h1f == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_31 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h20 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_32 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h21 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_33 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h22 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_34 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h23 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_35 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h24 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_36 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h25 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_37 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h26 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_38 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h27 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_39 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h28 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_40 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h29 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_41 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h2a == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_42 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h2b == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_43 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h2c == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_44 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h2d == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_45 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h2e == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_46 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h2f == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_47 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h30 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_48 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h31 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_49 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h32 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_50 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h33 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_51 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h34 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_52 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h35 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_53 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h36 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_54 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h37 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_55 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h38 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_56 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h39 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_57 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h3a == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_58 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h3b == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_59 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h3c == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_60 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h3d == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_61 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h3e == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_62 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h3f == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_63 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h40 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_64 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h41 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_65 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h42 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_66 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h43 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_67 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h44 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_68 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h45 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_69 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h46 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_70 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h47 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_71 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h48 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_72 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h49 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_73 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h4a == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_74 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h4b == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_75 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h4c == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_76 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h4d == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_77 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h4e == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_78 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h4f == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_79 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h50 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_80 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h51 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_81 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h52 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_82 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h53 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_83 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h54 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_84 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h55 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_85 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h56 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_86 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h57 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_87 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h58 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_88 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h59 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_89 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h5a == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_90 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h5b == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_91 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h5c == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_92 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h5d == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_93 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h5e == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_94 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h5f == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_95 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h60 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_96 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h61 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_97 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h62 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_98 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h63 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_99 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h64 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_100 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h65 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_101 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h66 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_102 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h67 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_103 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h68 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_104 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h69 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_105 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h6a == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_106 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h6b == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_107 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h6c == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_108 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h6d == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_109 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h6e == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_110 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h6f == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_111 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h70 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_112 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h71 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_113 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h72 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_114 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h73 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_115 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h74 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_116 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h75 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_117 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h76 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_118 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h77 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_119 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h78 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_120 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h79 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_121 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h7a == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_122 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h7b == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_123 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h7c == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_124 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h7d == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_125 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h7e == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_126 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h7f == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_127 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h80 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_128 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h81 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_129 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h82 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_130 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h83 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_131 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h84 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_132 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h85 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_133 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h86 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_134 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h87 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_135 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h88 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_136 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h89 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_137 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h8a == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_138 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h8b == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_139 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h8c == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_140 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h8d == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_141 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h8e == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_142 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h8f == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_143 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h90 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_144 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h91 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_145 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h92 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_146 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h93 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_147 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h94 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_148 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h95 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_149 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h96 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_150 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h97 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_151 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h98 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_152 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h99 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_153 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h9a == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_154 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h9b == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_155 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h9c == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_156 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h9d == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_157 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h9e == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_158 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h9f == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_159 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'ha0 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_160 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'ha1 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_161 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'ha2 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_162 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'ha3 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_163 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'ha4 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_164 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'ha5 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_165 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'ha6 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_166 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'ha7 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_167 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'ha8 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_168 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'ha9 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_169 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'haa == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_170 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'hab == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_171 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'hac == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_172 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'had == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_173 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'hae == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_174 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'haf == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_175 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'hb0 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_176 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'hb1 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_177 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'hb2 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_178 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'hb3 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_179 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'hb4 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_180 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'hb5 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_181 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'hb6 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_182 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'hb7 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_183 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'hb8 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_184 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'hb9 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_185 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'hba == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_186 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'hbb == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_187 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'hbc == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_188 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'hbd == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_189 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'hbe == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_190 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'hbf == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_191 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'hc0 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_192 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'hc1 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_193 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'hc2 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_194 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'hc3 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_195 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'hc4 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_196 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'hc5 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_197 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'hc6 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_198 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'hc7 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_199 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'hc8 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_200 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'hc9 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_201 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'hca == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_202 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'hcb == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_203 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'hcc == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_204 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'hcd == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_205 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'hce == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_206 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'hcf == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_207 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'hd0 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_208 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'hd1 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_209 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'hd2 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_210 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'hd3 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_211 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'hd4 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_212 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'hd5 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_213 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'hd6 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_214 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'hd7 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_215 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'hd8 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_216 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'hd9 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_217 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'hda == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_218 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'hdb == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_219 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'hdc == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_220 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'hdd == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_221 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'hde == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_222 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'hdf == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_223 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'he0 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_224 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'he1 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_225 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'he2 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_226 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'he3 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_227 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'he4 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_228 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'he5 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_229 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'he6 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_230 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'he7 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_231 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'he8 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_232 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'he9 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_233 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'hea == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_234 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'heb == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_235 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'hec == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_236 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'hed == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_237 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'hee == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_238 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'hef == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_239 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'hf0 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_240 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'hf1 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_241 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'hf2 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_242 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'hf3 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_243 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'hf4 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_244 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'hf5 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_245 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'hf6 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_246 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'hf7 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_247 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'hf8 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_248 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'hf9 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_249 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'hfa == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_250 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'hfb == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_251 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'hfc == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_252 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'hfd == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_253 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'hfe == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_254 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'hff == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_255 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h100 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_256 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h101 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_257 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h102 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_258 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h103 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_259 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h104 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_260 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h105 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_261 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h106 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_262 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h107 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_263 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h108 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_264 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h109 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_265 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h10a == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_266 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h10b == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_267 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h10c == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_268 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h10d == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_269 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h10e == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_270 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h10f == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_271 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h110 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_272 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h111 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_273 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h112 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_274 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h113 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_275 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h114 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_276 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h115 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_277 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h116 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_278 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h117 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_279 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h118 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_280 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h119 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_281 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h11a == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_282 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h11b == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_283 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h11c == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_284 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h11d == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_285 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h11e == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_286 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h11f == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_287 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h120 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_288 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h121 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_289 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h122 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_290 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h123 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_291 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h124 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_292 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h125 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_293 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h126 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_294 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h127 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_295 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h128 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_296 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h129 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_297 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h12a == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_298 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h12b == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_299 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h12c == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_300 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h12d == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_301 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h12e == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_302 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h12f == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_303 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h130 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_304 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h131 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_305 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h132 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_306 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h133 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_307 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h134 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_308 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h135 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_309 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h136 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_310 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h137 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_311 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h138 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_312 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h139 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_313 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h13a == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_314 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h13b == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_315 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h13c == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_316 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h13d == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_317 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h13e == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_318 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h13f == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_319 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h140 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_320 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h141 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_321 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h142 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_322 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h143 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_323 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h144 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_324 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h145 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_325 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h146 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_326 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h147 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_327 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h148 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_328 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h149 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_329 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h14a == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_330 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h14b == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_331 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h14c == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_332 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h14d == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_333 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h14e == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_334 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h14f == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_335 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h150 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_336 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h151 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_337 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h152 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_338 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h153 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_339 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h154 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_340 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h155 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_341 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h156 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_342 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h157 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_343 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h158 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_344 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h159 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_345 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h15a == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_346 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h15b == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_347 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h15c == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_348 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h15d == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_349 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h15e == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_350 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h15f == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_351 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h160 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_352 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h161 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_353 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h162 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_354 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h163 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_355 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h164 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_356 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h165 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_357 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h166 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_358 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h167 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_359 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h168 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_360 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h169 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_361 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h16a == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_362 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h16b == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_363 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h16c == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_364 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h16d == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_365 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h16e == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_366 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h16f == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_367 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h170 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_368 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h171 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_369 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h172 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_370 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h173 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_371 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h174 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_372 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h175 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_373 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h176 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_374 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h177 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_375 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h178 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_376 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h179 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_377 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h17a == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_378 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h17b == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_379 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h17c == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_380 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h17d == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_381 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h17e == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_382 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h17f == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_383 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h180 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_384 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h181 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_385 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h182 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_386 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h183 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_387 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h184 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_388 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h185 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_389 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h186 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_390 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h187 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_391 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h188 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_392 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h189 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_393 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h18a == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_394 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h18b == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_395 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h18c == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_396 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h18d == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_397 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h18e == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_398 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h18f == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_399 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h190 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_400 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h191 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_401 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h192 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_402 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h193 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_403 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h194 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_404 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h195 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_405 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h196 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_406 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h197 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_407 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h198 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_408 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h199 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_409 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h19a == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_410 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h19b == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_411 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h19c == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_412 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h19d == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_413 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h19e == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_414 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h19f == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_415 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h1a0 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_416 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h1a1 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_417 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h1a2 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_418 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h1a3 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_419 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h1a4 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_420 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h1a5 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_421 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h1a6 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_422 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h1a7 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_423 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h1a8 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_424 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h1a9 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_425 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h1aa == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_426 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h1ab == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_427 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h1ac == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_428 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h1ad == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_429 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h1ae == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_430 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h1af == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_431 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h1b0 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_432 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h1b1 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_433 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h1b2 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_434 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h1b3 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_435 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h1b4 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_436 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h1b5 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_437 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h1b6 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_438 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h1b7 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_439 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h1b8 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_440 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h1b9 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_441 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h1ba == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_442 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h1bb == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_443 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h1bc == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_444 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h1bd == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_445 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h1be == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_446 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h1bf == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_447 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h1c0 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_448 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h1c1 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_449 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h1c2 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_450 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h1c3 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_451 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h1c4 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_452 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h1c5 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_453 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h1c6 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_454 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h1c7 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_455 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h1c8 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_456 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h1c9 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_457 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h1ca == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_458 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h1cb == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_459 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h1cc == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_460 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h1cd == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_461 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h1ce == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_462 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h1cf == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_463 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h1d0 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_464 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h1d1 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_465 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h1d2 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_466 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h1d3 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_467 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h1d4 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_468 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h1d5 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_469 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h1d6 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_470 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h1d7 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_471 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h1d8 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_472 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h1d9 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_473 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h1da == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_474 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h1db == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_475 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h1dc == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_476 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h1dd == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_477 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h1de == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_478 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h1df == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_479 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h1e0 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_480 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h1e1 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_481 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h1e2 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_482 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h1e3 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_483 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h1e4 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_484 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h1e5 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_485 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h1e6 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_486 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h1e7 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_487 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h1e8 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_488 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h1e9 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_489 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h1ea == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_490 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h1eb == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_491 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h1ec == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_492 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h1ed == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_493 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h1ee == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_494 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h1ef == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_495 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h1f0 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_496 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h1f1 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_497 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h1f2 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_498 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h1f3 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_499 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h1f4 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_500 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h1f5 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_501 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h1f6 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_502 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h1f7 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_503 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h1f8 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_504 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h1f9 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_505 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h1fa == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_506 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h1fb == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_507 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h1fc == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_508 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h1fd == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_509 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h1fe == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_510 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h1ff == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_511 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h200 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_512 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h201 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_513 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h202 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_514 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h203 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_515 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h204 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_516 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h205 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_517 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h206 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_518 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h207 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_519 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h208 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_520 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h209 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_521 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h20a == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_522 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h20b == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_523 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h20c == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_524 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h20d == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_525 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h20e == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_526 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h20f == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_527 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h210 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_528 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h211 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_529 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h212 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_530 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h213 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_531 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h214 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_532 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h215 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_533 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h216 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_534 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h217 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_535 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h218 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_536 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h219 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_537 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h21a == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_538 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h21b == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_539 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h21c == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_540 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h21d == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_541 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h21e == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_542 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h21f == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_543 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h220 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_544 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h221 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_545 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h222 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_546 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h223 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_547 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h224 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_548 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h225 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_549 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h226 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_550 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h227 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_551 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h228 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_552 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h229 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_553 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h22a == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_554 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h22b == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_555 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h22c == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_556 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h22d == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_557 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h22e == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_558 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h22f == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_559 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h230 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_560 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h231 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_561 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h232 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_562 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h233 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_563 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h234 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_564 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h235 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_565 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h236 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_566 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h237 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_567 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h238 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_568 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h239 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_569 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h23a == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_570 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h23b == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_571 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h23c == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_572 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h23d == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_573 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h23e == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_574 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h23f == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_575 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h240 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_576 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h241 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_577 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h242 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_578 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h243 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_579 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h244 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_580 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h245 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_581 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h246 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_582 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h247 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_583 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h248 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_584 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h249 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_585 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h24a == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_586 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h24b == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_587 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h24c == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_588 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h24d == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_589 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h24e == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_590 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h24f == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_591 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h250 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_592 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h251 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_593 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h252 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_594 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h253 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_595 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h254 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_596 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h255 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_597 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h256 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_598 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h257 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_599 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h258 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_600 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h259 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_601 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h25a == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_602 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h25b == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_603 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h25c == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_604 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h25d == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_605 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h25e == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_606 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h25f == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_607 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h260 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_608 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h261 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_609 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h262 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_610 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h263 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_611 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h264 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_612 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h265 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_613 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h266 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_614 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h267 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_615 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h268 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_616 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h269 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_617 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h26a == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_618 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h26b == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_619 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h26c == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_620 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h26d == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_621 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h26e == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_622 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h26f == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_623 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h270 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_624 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h271 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_625 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h272 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_626 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h273 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_627 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h274 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_628 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h275 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_629 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h276 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_630 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h277 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_631 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h278 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_632 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h279 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_633 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h27a == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_634 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h27b == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_635 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h27c == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_636 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h27d == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_637 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h27e == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_638 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h27f == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_639 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h280 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_640 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h281 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_641 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h282 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_642 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h283 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_643 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h284 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_644 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h285 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_645 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h286 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_646 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h287 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_647 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h288 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_648 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h289 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_649 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h28a == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_650 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h28b == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_651 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h28c == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_652 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h28d == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_653 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h28e == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_654 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h28f == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_655 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h290 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_656 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h291 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_657 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h292 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_658 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h293 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_659 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h294 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_660 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h295 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_661 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h296 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_662 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h297 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_663 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h298 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_664 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h299 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_665 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h29a == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_666 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h29b == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_667 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h29c == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_668 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h29d == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_669 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h29e == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_670 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h29f == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_671 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h2a0 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_672 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h2a1 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_673 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h2a2 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_674 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h2a3 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_675 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h2a4 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_676 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h2a5 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_677 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h2a6 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_678 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h2a7 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_679 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h2a8 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_680 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h2a9 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_681 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h2aa == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_682 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h2ab == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_683 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h2ac == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_684 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h2ad == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_685 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h2ae == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_686 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h2af == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_687 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h2b0 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_688 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h2b1 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_689 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h2b2 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_690 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h2b3 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_691 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h2b4 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_692 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h2b5 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_693 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h2b6 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_694 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h2b7 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_695 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h2b8 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_696 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h2b9 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_697 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h2ba == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_698 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h2bb == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_699 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h2bc == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_700 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h2bd == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_701 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h2be == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_702 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h2bf == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_703 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h2c0 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_704 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h2c1 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_705 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h2c2 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_706 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h2c3 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_707 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h2c4 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_708 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h2c5 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_709 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h2c6 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_710 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h2c7 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_711 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h2c8 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_712 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h2c9 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_713 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h2ca == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_714 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h2cb == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_715 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h2cc == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_716 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h2cd == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_717 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h2ce == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_718 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h2cf == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_719 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h2d0 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_720 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h2d1 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_721 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h2d2 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_722 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h2d3 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_723 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h2d4 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_724 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h2d5 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_725 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h2d6 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_726 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h2d7 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_727 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h2d8 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_728 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h2d9 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_729 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h2da == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_730 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h2db == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_731 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h2dc == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_732 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h2dd == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_733 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h2de == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_734 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h2df == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_735 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h2e0 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_736 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h2e1 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_737 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h2e2 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_738 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h2e3 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_739 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h2e4 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_740 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h2e5 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_741 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h2e6 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_742 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h2e7 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_743 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h2e8 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_744 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h2e9 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_745 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h2ea == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_746 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h2eb == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_747 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h2ec == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_748 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h2ed == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_749 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h2ee == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_750 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h2ef == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_751 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h2f0 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_752 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h2f1 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_753 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h2f2 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_754 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h2f3 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_755 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h2f4 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_756 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h2f5 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_757 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h2f6 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_758 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h2f7 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_759 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h2f8 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_760 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h2f9 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_761 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h2fa == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_762 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h2fb == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_763 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h2fc == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_764 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h2fd == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_765 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h2fe == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_766 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h2ff == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_767 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h300 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_768 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h301 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_769 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h302 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_770 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h303 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_771 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h304 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_772 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h305 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_773 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h306 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_774 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h307 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_775 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h308 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_776 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h309 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_777 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h30a == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_778 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h30b == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_779 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h30c == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_780 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h30d == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_781 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h30e == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_782 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h30f == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_783 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h310 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_784 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h311 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_785 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h312 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_786 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h313 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_787 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h314 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_788 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h315 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_789 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h316 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_790 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h317 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_791 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h318 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_792 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h319 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_793 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h31a == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_794 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h31b == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_795 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h31c == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_796 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h31d == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_797 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h31e == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_798 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h31f == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_799 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h320 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_800 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h321 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_801 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h322 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_802 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h323 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_803 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h324 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_804 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h325 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_805 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h326 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_806 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h327 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_807 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h328 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_808 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h329 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_809 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h32a == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_810 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h32b == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_811 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h32c == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_812 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h32d == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_813 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h32e == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_814 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h32f == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_815 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h330 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_816 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h331 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_817 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h332 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_818 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h333 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_819 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h334 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_820 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h335 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_821 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h336 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_822 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h337 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_823 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h338 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_824 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h339 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_825 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h33a == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_826 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h33b == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_827 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h33c == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_828 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h33d == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_829 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h33e == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_830 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h33f == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_831 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h340 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_832 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h341 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_833 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h342 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_834 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h343 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_835 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h344 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_836 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h345 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_837 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h346 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_838 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h347 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_839 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h348 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_840 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h349 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_841 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h34a == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_842 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h34b == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_843 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h34c == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_844 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h34d == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_845 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h34e == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_846 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h34f == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_847 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h350 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_848 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h351 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_849 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h352 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_850 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h353 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_851 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h354 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_852 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h355 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_853 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h356 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_854 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h357 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_855 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h358 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_856 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h359 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_857 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h35a == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_858 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h35b == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_859 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h35c == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_860 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h35d == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_861 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h35e == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_862 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h35f == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_863 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h360 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_864 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h361 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_865 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h362 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_866 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h363 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_867 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h364 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_868 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h365 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_869 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h366 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_870 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h367 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_871 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h368 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_872 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h369 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_873 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h36a == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_874 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h36b == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_875 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h36c == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_876 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h36d == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_877 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h36e == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_878 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h36f == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_879 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h370 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_880 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h371 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_881 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h372 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_882 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h373 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_883 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h374 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_884 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h375 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_885 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h376 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_886 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h377 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_887 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h378 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_888 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h379 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_889 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h37a == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_890 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h37b == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_891 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h37c == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_892 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h37d == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_893 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h37e == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_894 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h37f == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_895 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h380 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_896 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h381 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_897 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h382 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_898 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h383 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_899 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h384 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_900 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h385 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_901 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h386 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_902 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h387 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_903 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h388 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_904 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h389 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_905 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h38a == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_906 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h38b == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_907 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h38c == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_908 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h38d == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_909 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h38e == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_910 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h38f == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_911 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h390 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_912 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h391 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_913 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h392 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_914 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h393 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_915 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h394 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_916 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h395 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_917 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h396 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_918 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h397 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_919 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h398 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_920 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h399 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_921 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h39a == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_922 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h39b == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_923 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h39c == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_924 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h39d == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_925 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h39e == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_926 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h39f == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_927 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h3a0 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_928 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h3a1 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_929 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h3a2 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_930 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h3a3 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_931 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h3a4 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_932 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h3a5 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_933 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h3a6 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_934 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h3a7 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_935 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h3a8 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_936 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h3a9 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_937 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h3aa == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_938 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h3ab == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_939 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h3ac == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_940 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h3ad == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_941 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h3ae == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_942 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h3af == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_943 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h3b0 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_944 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h3b1 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_945 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h3b2 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_946 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h3b3 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_947 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h3b4 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_948 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h3b5 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_949 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h3b6 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_950 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h3b7 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_951 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h3b8 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_952 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h3b9 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_953 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h3ba == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_954 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h3bb == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_955 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h3bc == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_956 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h3bd == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_957 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h3be == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_958 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h3bf == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_959 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h3c0 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_960 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h3c1 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_961 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h3c2 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_962 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h3c3 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_963 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h3c4 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_964 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h3c5 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_965 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h3c6 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_966 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h3c7 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_967 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h3c8 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_968 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h3c9 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_969 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h3ca == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_970 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h3cb == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_971 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h3cc == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_972 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h3cd == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_973 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h3ce == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_974 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h3cf == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_975 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h3d0 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_976 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h3d1 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_977 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h3d2 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_978 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h3d3 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_979 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h3d4 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_980 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h3d5 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_981 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h3d6 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_982 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h3d7 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_983 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h3d8 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_984 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h3d9 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_985 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h3da == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_986 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h3db == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_987 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h3dc == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_988 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h3dd == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_989 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h3de == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_990 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h3df == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_991 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h3e0 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_992 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h3e1 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_993 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h3e2 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_994 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h3e3 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_995 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h3e4 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_996 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h3e5 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_997 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h3e6 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_998 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h3e7 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_999 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h3e8 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_1000 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h3e9 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_1001 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h3ea == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_1002 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h3eb == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_1003 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h3ec == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_1004 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h3ed == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_1005 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h3ee == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_1006 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h3ef == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_1007 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h3f0 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_1008 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h3f1 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_1009 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h3f2 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_1010 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h3f3 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_1011 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h3f4 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_1012 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h3f5 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_1013 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h3f6 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_1014 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h3f7 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_1015 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h3f8 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_1016 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h3f9 == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_1017 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h3fa == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_1018 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h3fb == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_1019 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h3fc == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_1020 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h3fd == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_1021 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h3fe == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_1022 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
    if (_T_2) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 42:62]
      if (10'h3ff == WritePtr[9:0]) begin // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
        FifoCell_1023 <= io_Writer_WriteData; // @[src/main/scala/fifo_pkg/FifoPkg.scala 43:43]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  WritePtr = _RAND_0[10:0];
  _RAND_1 = {1{`RANDOM}};
  ReadPtr = _RAND_1[10:0];
  _RAND_2 = {1{`RANDOM}};
  FifoCell_0 = _RAND_2[8:0];
  _RAND_3 = {1{`RANDOM}};
  FifoCell_1 = _RAND_3[8:0];
  _RAND_4 = {1{`RANDOM}};
  FifoCell_2 = _RAND_4[8:0];
  _RAND_5 = {1{`RANDOM}};
  FifoCell_3 = _RAND_5[8:0];
  _RAND_6 = {1{`RANDOM}};
  FifoCell_4 = _RAND_6[8:0];
  _RAND_7 = {1{`RANDOM}};
  FifoCell_5 = _RAND_7[8:0];
  _RAND_8 = {1{`RANDOM}};
  FifoCell_6 = _RAND_8[8:0];
  _RAND_9 = {1{`RANDOM}};
  FifoCell_7 = _RAND_9[8:0];
  _RAND_10 = {1{`RANDOM}};
  FifoCell_8 = _RAND_10[8:0];
  _RAND_11 = {1{`RANDOM}};
  FifoCell_9 = _RAND_11[8:0];
  _RAND_12 = {1{`RANDOM}};
  FifoCell_10 = _RAND_12[8:0];
  _RAND_13 = {1{`RANDOM}};
  FifoCell_11 = _RAND_13[8:0];
  _RAND_14 = {1{`RANDOM}};
  FifoCell_12 = _RAND_14[8:0];
  _RAND_15 = {1{`RANDOM}};
  FifoCell_13 = _RAND_15[8:0];
  _RAND_16 = {1{`RANDOM}};
  FifoCell_14 = _RAND_16[8:0];
  _RAND_17 = {1{`RANDOM}};
  FifoCell_15 = _RAND_17[8:0];
  _RAND_18 = {1{`RANDOM}};
  FifoCell_16 = _RAND_18[8:0];
  _RAND_19 = {1{`RANDOM}};
  FifoCell_17 = _RAND_19[8:0];
  _RAND_20 = {1{`RANDOM}};
  FifoCell_18 = _RAND_20[8:0];
  _RAND_21 = {1{`RANDOM}};
  FifoCell_19 = _RAND_21[8:0];
  _RAND_22 = {1{`RANDOM}};
  FifoCell_20 = _RAND_22[8:0];
  _RAND_23 = {1{`RANDOM}};
  FifoCell_21 = _RAND_23[8:0];
  _RAND_24 = {1{`RANDOM}};
  FifoCell_22 = _RAND_24[8:0];
  _RAND_25 = {1{`RANDOM}};
  FifoCell_23 = _RAND_25[8:0];
  _RAND_26 = {1{`RANDOM}};
  FifoCell_24 = _RAND_26[8:0];
  _RAND_27 = {1{`RANDOM}};
  FifoCell_25 = _RAND_27[8:0];
  _RAND_28 = {1{`RANDOM}};
  FifoCell_26 = _RAND_28[8:0];
  _RAND_29 = {1{`RANDOM}};
  FifoCell_27 = _RAND_29[8:0];
  _RAND_30 = {1{`RANDOM}};
  FifoCell_28 = _RAND_30[8:0];
  _RAND_31 = {1{`RANDOM}};
  FifoCell_29 = _RAND_31[8:0];
  _RAND_32 = {1{`RANDOM}};
  FifoCell_30 = _RAND_32[8:0];
  _RAND_33 = {1{`RANDOM}};
  FifoCell_31 = _RAND_33[8:0];
  _RAND_34 = {1{`RANDOM}};
  FifoCell_32 = _RAND_34[8:0];
  _RAND_35 = {1{`RANDOM}};
  FifoCell_33 = _RAND_35[8:0];
  _RAND_36 = {1{`RANDOM}};
  FifoCell_34 = _RAND_36[8:0];
  _RAND_37 = {1{`RANDOM}};
  FifoCell_35 = _RAND_37[8:0];
  _RAND_38 = {1{`RANDOM}};
  FifoCell_36 = _RAND_38[8:0];
  _RAND_39 = {1{`RANDOM}};
  FifoCell_37 = _RAND_39[8:0];
  _RAND_40 = {1{`RANDOM}};
  FifoCell_38 = _RAND_40[8:0];
  _RAND_41 = {1{`RANDOM}};
  FifoCell_39 = _RAND_41[8:0];
  _RAND_42 = {1{`RANDOM}};
  FifoCell_40 = _RAND_42[8:0];
  _RAND_43 = {1{`RANDOM}};
  FifoCell_41 = _RAND_43[8:0];
  _RAND_44 = {1{`RANDOM}};
  FifoCell_42 = _RAND_44[8:0];
  _RAND_45 = {1{`RANDOM}};
  FifoCell_43 = _RAND_45[8:0];
  _RAND_46 = {1{`RANDOM}};
  FifoCell_44 = _RAND_46[8:0];
  _RAND_47 = {1{`RANDOM}};
  FifoCell_45 = _RAND_47[8:0];
  _RAND_48 = {1{`RANDOM}};
  FifoCell_46 = _RAND_48[8:0];
  _RAND_49 = {1{`RANDOM}};
  FifoCell_47 = _RAND_49[8:0];
  _RAND_50 = {1{`RANDOM}};
  FifoCell_48 = _RAND_50[8:0];
  _RAND_51 = {1{`RANDOM}};
  FifoCell_49 = _RAND_51[8:0];
  _RAND_52 = {1{`RANDOM}};
  FifoCell_50 = _RAND_52[8:0];
  _RAND_53 = {1{`RANDOM}};
  FifoCell_51 = _RAND_53[8:0];
  _RAND_54 = {1{`RANDOM}};
  FifoCell_52 = _RAND_54[8:0];
  _RAND_55 = {1{`RANDOM}};
  FifoCell_53 = _RAND_55[8:0];
  _RAND_56 = {1{`RANDOM}};
  FifoCell_54 = _RAND_56[8:0];
  _RAND_57 = {1{`RANDOM}};
  FifoCell_55 = _RAND_57[8:0];
  _RAND_58 = {1{`RANDOM}};
  FifoCell_56 = _RAND_58[8:0];
  _RAND_59 = {1{`RANDOM}};
  FifoCell_57 = _RAND_59[8:0];
  _RAND_60 = {1{`RANDOM}};
  FifoCell_58 = _RAND_60[8:0];
  _RAND_61 = {1{`RANDOM}};
  FifoCell_59 = _RAND_61[8:0];
  _RAND_62 = {1{`RANDOM}};
  FifoCell_60 = _RAND_62[8:0];
  _RAND_63 = {1{`RANDOM}};
  FifoCell_61 = _RAND_63[8:0];
  _RAND_64 = {1{`RANDOM}};
  FifoCell_62 = _RAND_64[8:0];
  _RAND_65 = {1{`RANDOM}};
  FifoCell_63 = _RAND_65[8:0];
  _RAND_66 = {1{`RANDOM}};
  FifoCell_64 = _RAND_66[8:0];
  _RAND_67 = {1{`RANDOM}};
  FifoCell_65 = _RAND_67[8:0];
  _RAND_68 = {1{`RANDOM}};
  FifoCell_66 = _RAND_68[8:0];
  _RAND_69 = {1{`RANDOM}};
  FifoCell_67 = _RAND_69[8:0];
  _RAND_70 = {1{`RANDOM}};
  FifoCell_68 = _RAND_70[8:0];
  _RAND_71 = {1{`RANDOM}};
  FifoCell_69 = _RAND_71[8:0];
  _RAND_72 = {1{`RANDOM}};
  FifoCell_70 = _RAND_72[8:0];
  _RAND_73 = {1{`RANDOM}};
  FifoCell_71 = _RAND_73[8:0];
  _RAND_74 = {1{`RANDOM}};
  FifoCell_72 = _RAND_74[8:0];
  _RAND_75 = {1{`RANDOM}};
  FifoCell_73 = _RAND_75[8:0];
  _RAND_76 = {1{`RANDOM}};
  FifoCell_74 = _RAND_76[8:0];
  _RAND_77 = {1{`RANDOM}};
  FifoCell_75 = _RAND_77[8:0];
  _RAND_78 = {1{`RANDOM}};
  FifoCell_76 = _RAND_78[8:0];
  _RAND_79 = {1{`RANDOM}};
  FifoCell_77 = _RAND_79[8:0];
  _RAND_80 = {1{`RANDOM}};
  FifoCell_78 = _RAND_80[8:0];
  _RAND_81 = {1{`RANDOM}};
  FifoCell_79 = _RAND_81[8:0];
  _RAND_82 = {1{`RANDOM}};
  FifoCell_80 = _RAND_82[8:0];
  _RAND_83 = {1{`RANDOM}};
  FifoCell_81 = _RAND_83[8:0];
  _RAND_84 = {1{`RANDOM}};
  FifoCell_82 = _RAND_84[8:0];
  _RAND_85 = {1{`RANDOM}};
  FifoCell_83 = _RAND_85[8:0];
  _RAND_86 = {1{`RANDOM}};
  FifoCell_84 = _RAND_86[8:0];
  _RAND_87 = {1{`RANDOM}};
  FifoCell_85 = _RAND_87[8:0];
  _RAND_88 = {1{`RANDOM}};
  FifoCell_86 = _RAND_88[8:0];
  _RAND_89 = {1{`RANDOM}};
  FifoCell_87 = _RAND_89[8:0];
  _RAND_90 = {1{`RANDOM}};
  FifoCell_88 = _RAND_90[8:0];
  _RAND_91 = {1{`RANDOM}};
  FifoCell_89 = _RAND_91[8:0];
  _RAND_92 = {1{`RANDOM}};
  FifoCell_90 = _RAND_92[8:0];
  _RAND_93 = {1{`RANDOM}};
  FifoCell_91 = _RAND_93[8:0];
  _RAND_94 = {1{`RANDOM}};
  FifoCell_92 = _RAND_94[8:0];
  _RAND_95 = {1{`RANDOM}};
  FifoCell_93 = _RAND_95[8:0];
  _RAND_96 = {1{`RANDOM}};
  FifoCell_94 = _RAND_96[8:0];
  _RAND_97 = {1{`RANDOM}};
  FifoCell_95 = _RAND_97[8:0];
  _RAND_98 = {1{`RANDOM}};
  FifoCell_96 = _RAND_98[8:0];
  _RAND_99 = {1{`RANDOM}};
  FifoCell_97 = _RAND_99[8:0];
  _RAND_100 = {1{`RANDOM}};
  FifoCell_98 = _RAND_100[8:0];
  _RAND_101 = {1{`RANDOM}};
  FifoCell_99 = _RAND_101[8:0];
  _RAND_102 = {1{`RANDOM}};
  FifoCell_100 = _RAND_102[8:0];
  _RAND_103 = {1{`RANDOM}};
  FifoCell_101 = _RAND_103[8:0];
  _RAND_104 = {1{`RANDOM}};
  FifoCell_102 = _RAND_104[8:0];
  _RAND_105 = {1{`RANDOM}};
  FifoCell_103 = _RAND_105[8:0];
  _RAND_106 = {1{`RANDOM}};
  FifoCell_104 = _RAND_106[8:0];
  _RAND_107 = {1{`RANDOM}};
  FifoCell_105 = _RAND_107[8:0];
  _RAND_108 = {1{`RANDOM}};
  FifoCell_106 = _RAND_108[8:0];
  _RAND_109 = {1{`RANDOM}};
  FifoCell_107 = _RAND_109[8:0];
  _RAND_110 = {1{`RANDOM}};
  FifoCell_108 = _RAND_110[8:0];
  _RAND_111 = {1{`RANDOM}};
  FifoCell_109 = _RAND_111[8:0];
  _RAND_112 = {1{`RANDOM}};
  FifoCell_110 = _RAND_112[8:0];
  _RAND_113 = {1{`RANDOM}};
  FifoCell_111 = _RAND_113[8:0];
  _RAND_114 = {1{`RANDOM}};
  FifoCell_112 = _RAND_114[8:0];
  _RAND_115 = {1{`RANDOM}};
  FifoCell_113 = _RAND_115[8:0];
  _RAND_116 = {1{`RANDOM}};
  FifoCell_114 = _RAND_116[8:0];
  _RAND_117 = {1{`RANDOM}};
  FifoCell_115 = _RAND_117[8:0];
  _RAND_118 = {1{`RANDOM}};
  FifoCell_116 = _RAND_118[8:0];
  _RAND_119 = {1{`RANDOM}};
  FifoCell_117 = _RAND_119[8:0];
  _RAND_120 = {1{`RANDOM}};
  FifoCell_118 = _RAND_120[8:0];
  _RAND_121 = {1{`RANDOM}};
  FifoCell_119 = _RAND_121[8:0];
  _RAND_122 = {1{`RANDOM}};
  FifoCell_120 = _RAND_122[8:0];
  _RAND_123 = {1{`RANDOM}};
  FifoCell_121 = _RAND_123[8:0];
  _RAND_124 = {1{`RANDOM}};
  FifoCell_122 = _RAND_124[8:0];
  _RAND_125 = {1{`RANDOM}};
  FifoCell_123 = _RAND_125[8:0];
  _RAND_126 = {1{`RANDOM}};
  FifoCell_124 = _RAND_126[8:0];
  _RAND_127 = {1{`RANDOM}};
  FifoCell_125 = _RAND_127[8:0];
  _RAND_128 = {1{`RANDOM}};
  FifoCell_126 = _RAND_128[8:0];
  _RAND_129 = {1{`RANDOM}};
  FifoCell_127 = _RAND_129[8:0];
  _RAND_130 = {1{`RANDOM}};
  FifoCell_128 = _RAND_130[8:0];
  _RAND_131 = {1{`RANDOM}};
  FifoCell_129 = _RAND_131[8:0];
  _RAND_132 = {1{`RANDOM}};
  FifoCell_130 = _RAND_132[8:0];
  _RAND_133 = {1{`RANDOM}};
  FifoCell_131 = _RAND_133[8:0];
  _RAND_134 = {1{`RANDOM}};
  FifoCell_132 = _RAND_134[8:0];
  _RAND_135 = {1{`RANDOM}};
  FifoCell_133 = _RAND_135[8:0];
  _RAND_136 = {1{`RANDOM}};
  FifoCell_134 = _RAND_136[8:0];
  _RAND_137 = {1{`RANDOM}};
  FifoCell_135 = _RAND_137[8:0];
  _RAND_138 = {1{`RANDOM}};
  FifoCell_136 = _RAND_138[8:0];
  _RAND_139 = {1{`RANDOM}};
  FifoCell_137 = _RAND_139[8:0];
  _RAND_140 = {1{`RANDOM}};
  FifoCell_138 = _RAND_140[8:0];
  _RAND_141 = {1{`RANDOM}};
  FifoCell_139 = _RAND_141[8:0];
  _RAND_142 = {1{`RANDOM}};
  FifoCell_140 = _RAND_142[8:0];
  _RAND_143 = {1{`RANDOM}};
  FifoCell_141 = _RAND_143[8:0];
  _RAND_144 = {1{`RANDOM}};
  FifoCell_142 = _RAND_144[8:0];
  _RAND_145 = {1{`RANDOM}};
  FifoCell_143 = _RAND_145[8:0];
  _RAND_146 = {1{`RANDOM}};
  FifoCell_144 = _RAND_146[8:0];
  _RAND_147 = {1{`RANDOM}};
  FifoCell_145 = _RAND_147[8:0];
  _RAND_148 = {1{`RANDOM}};
  FifoCell_146 = _RAND_148[8:0];
  _RAND_149 = {1{`RANDOM}};
  FifoCell_147 = _RAND_149[8:0];
  _RAND_150 = {1{`RANDOM}};
  FifoCell_148 = _RAND_150[8:0];
  _RAND_151 = {1{`RANDOM}};
  FifoCell_149 = _RAND_151[8:0];
  _RAND_152 = {1{`RANDOM}};
  FifoCell_150 = _RAND_152[8:0];
  _RAND_153 = {1{`RANDOM}};
  FifoCell_151 = _RAND_153[8:0];
  _RAND_154 = {1{`RANDOM}};
  FifoCell_152 = _RAND_154[8:0];
  _RAND_155 = {1{`RANDOM}};
  FifoCell_153 = _RAND_155[8:0];
  _RAND_156 = {1{`RANDOM}};
  FifoCell_154 = _RAND_156[8:0];
  _RAND_157 = {1{`RANDOM}};
  FifoCell_155 = _RAND_157[8:0];
  _RAND_158 = {1{`RANDOM}};
  FifoCell_156 = _RAND_158[8:0];
  _RAND_159 = {1{`RANDOM}};
  FifoCell_157 = _RAND_159[8:0];
  _RAND_160 = {1{`RANDOM}};
  FifoCell_158 = _RAND_160[8:0];
  _RAND_161 = {1{`RANDOM}};
  FifoCell_159 = _RAND_161[8:0];
  _RAND_162 = {1{`RANDOM}};
  FifoCell_160 = _RAND_162[8:0];
  _RAND_163 = {1{`RANDOM}};
  FifoCell_161 = _RAND_163[8:0];
  _RAND_164 = {1{`RANDOM}};
  FifoCell_162 = _RAND_164[8:0];
  _RAND_165 = {1{`RANDOM}};
  FifoCell_163 = _RAND_165[8:0];
  _RAND_166 = {1{`RANDOM}};
  FifoCell_164 = _RAND_166[8:0];
  _RAND_167 = {1{`RANDOM}};
  FifoCell_165 = _RAND_167[8:0];
  _RAND_168 = {1{`RANDOM}};
  FifoCell_166 = _RAND_168[8:0];
  _RAND_169 = {1{`RANDOM}};
  FifoCell_167 = _RAND_169[8:0];
  _RAND_170 = {1{`RANDOM}};
  FifoCell_168 = _RAND_170[8:0];
  _RAND_171 = {1{`RANDOM}};
  FifoCell_169 = _RAND_171[8:0];
  _RAND_172 = {1{`RANDOM}};
  FifoCell_170 = _RAND_172[8:0];
  _RAND_173 = {1{`RANDOM}};
  FifoCell_171 = _RAND_173[8:0];
  _RAND_174 = {1{`RANDOM}};
  FifoCell_172 = _RAND_174[8:0];
  _RAND_175 = {1{`RANDOM}};
  FifoCell_173 = _RAND_175[8:0];
  _RAND_176 = {1{`RANDOM}};
  FifoCell_174 = _RAND_176[8:0];
  _RAND_177 = {1{`RANDOM}};
  FifoCell_175 = _RAND_177[8:0];
  _RAND_178 = {1{`RANDOM}};
  FifoCell_176 = _RAND_178[8:0];
  _RAND_179 = {1{`RANDOM}};
  FifoCell_177 = _RAND_179[8:0];
  _RAND_180 = {1{`RANDOM}};
  FifoCell_178 = _RAND_180[8:0];
  _RAND_181 = {1{`RANDOM}};
  FifoCell_179 = _RAND_181[8:0];
  _RAND_182 = {1{`RANDOM}};
  FifoCell_180 = _RAND_182[8:0];
  _RAND_183 = {1{`RANDOM}};
  FifoCell_181 = _RAND_183[8:0];
  _RAND_184 = {1{`RANDOM}};
  FifoCell_182 = _RAND_184[8:0];
  _RAND_185 = {1{`RANDOM}};
  FifoCell_183 = _RAND_185[8:0];
  _RAND_186 = {1{`RANDOM}};
  FifoCell_184 = _RAND_186[8:0];
  _RAND_187 = {1{`RANDOM}};
  FifoCell_185 = _RAND_187[8:0];
  _RAND_188 = {1{`RANDOM}};
  FifoCell_186 = _RAND_188[8:0];
  _RAND_189 = {1{`RANDOM}};
  FifoCell_187 = _RAND_189[8:0];
  _RAND_190 = {1{`RANDOM}};
  FifoCell_188 = _RAND_190[8:0];
  _RAND_191 = {1{`RANDOM}};
  FifoCell_189 = _RAND_191[8:0];
  _RAND_192 = {1{`RANDOM}};
  FifoCell_190 = _RAND_192[8:0];
  _RAND_193 = {1{`RANDOM}};
  FifoCell_191 = _RAND_193[8:0];
  _RAND_194 = {1{`RANDOM}};
  FifoCell_192 = _RAND_194[8:0];
  _RAND_195 = {1{`RANDOM}};
  FifoCell_193 = _RAND_195[8:0];
  _RAND_196 = {1{`RANDOM}};
  FifoCell_194 = _RAND_196[8:0];
  _RAND_197 = {1{`RANDOM}};
  FifoCell_195 = _RAND_197[8:0];
  _RAND_198 = {1{`RANDOM}};
  FifoCell_196 = _RAND_198[8:0];
  _RAND_199 = {1{`RANDOM}};
  FifoCell_197 = _RAND_199[8:0];
  _RAND_200 = {1{`RANDOM}};
  FifoCell_198 = _RAND_200[8:0];
  _RAND_201 = {1{`RANDOM}};
  FifoCell_199 = _RAND_201[8:0];
  _RAND_202 = {1{`RANDOM}};
  FifoCell_200 = _RAND_202[8:0];
  _RAND_203 = {1{`RANDOM}};
  FifoCell_201 = _RAND_203[8:0];
  _RAND_204 = {1{`RANDOM}};
  FifoCell_202 = _RAND_204[8:0];
  _RAND_205 = {1{`RANDOM}};
  FifoCell_203 = _RAND_205[8:0];
  _RAND_206 = {1{`RANDOM}};
  FifoCell_204 = _RAND_206[8:0];
  _RAND_207 = {1{`RANDOM}};
  FifoCell_205 = _RAND_207[8:0];
  _RAND_208 = {1{`RANDOM}};
  FifoCell_206 = _RAND_208[8:0];
  _RAND_209 = {1{`RANDOM}};
  FifoCell_207 = _RAND_209[8:0];
  _RAND_210 = {1{`RANDOM}};
  FifoCell_208 = _RAND_210[8:0];
  _RAND_211 = {1{`RANDOM}};
  FifoCell_209 = _RAND_211[8:0];
  _RAND_212 = {1{`RANDOM}};
  FifoCell_210 = _RAND_212[8:0];
  _RAND_213 = {1{`RANDOM}};
  FifoCell_211 = _RAND_213[8:0];
  _RAND_214 = {1{`RANDOM}};
  FifoCell_212 = _RAND_214[8:0];
  _RAND_215 = {1{`RANDOM}};
  FifoCell_213 = _RAND_215[8:0];
  _RAND_216 = {1{`RANDOM}};
  FifoCell_214 = _RAND_216[8:0];
  _RAND_217 = {1{`RANDOM}};
  FifoCell_215 = _RAND_217[8:0];
  _RAND_218 = {1{`RANDOM}};
  FifoCell_216 = _RAND_218[8:0];
  _RAND_219 = {1{`RANDOM}};
  FifoCell_217 = _RAND_219[8:0];
  _RAND_220 = {1{`RANDOM}};
  FifoCell_218 = _RAND_220[8:0];
  _RAND_221 = {1{`RANDOM}};
  FifoCell_219 = _RAND_221[8:0];
  _RAND_222 = {1{`RANDOM}};
  FifoCell_220 = _RAND_222[8:0];
  _RAND_223 = {1{`RANDOM}};
  FifoCell_221 = _RAND_223[8:0];
  _RAND_224 = {1{`RANDOM}};
  FifoCell_222 = _RAND_224[8:0];
  _RAND_225 = {1{`RANDOM}};
  FifoCell_223 = _RAND_225[8:0];
  _RAND_226 = {1{`RANDOM}};
  FifoCell_224 = _RAND_226[8:0];
  _RAND_227 = {1{`RANDOM}};
  FifoCell_225 = _RAND_227[8:0];
  _RAND_228 = {1{`RANDOM}};
  FifoCell_226 = _RAND_228[8:0];
  _RAND_229 = {1{`RANDOM}};
  FifoCell_227 = _RAND_229[8:0];
  _RAND_230 = {1{`RANDOM}};
  FifoCell_228 = _RAND_230[8:0];
  _RAND_231 = {1{`RANDOM}};
  FifoCell_229 = _RAND_231[8:0];
  _RAND_232 = {1{`RANDOM}};
  FifoCell_230 = _RAND_232[8:0];
  _RAND_233 = {1{`RANDOM}};
  FifoCell_231 = _RAND_233[8:0];
  _RAND_234 = {1{`RANDOM}};
  FifoCell_232 = _RAND_234[8:0];
  _RAND_235 = {1{`RANDOM}};
  FifoCell_233 = _RAND_235[8:0];
  _RAND_236 = {1{`RANDOM}};
  FifoCell_234 = _RAND_236[8:0];
  _RAND_237 = {1{`RANDOM}};
  FifoCell_235 = _RAND_237[8:0];
  _RAND_238 = {1{`RANDOM}};
  FifoCell_236 = _RAND_238[8:0];
  _RAND_239 = {1{`RANDOM}};
  FifoCell_237 = _RAND_239[8:0];
  _RAND_240 = {1{`RANDOM}};
  FifoCell_238 = _RAND_240[8:0];
  _RAND_241 = {1{`RANDOM}};
  FifoCell_239 = _RAND_241[8:0];
  _RAND_242 = {1{`RANDOM}};
  FifoCell_240 = _RAND_242[8:0];
  _RAND_243 = {1{`RANDOM}};
  FifoCell_241 = _RAND_243[8:0];
  _RAND_244 = {1{`RANDOM}};
  FifoCell_242 = _RAND_244[8:0];
  _RAND_245 = {1{`RANDOM}};
  FifoCell_243 = _RAND_245[8:0];
  _RAND_246 = {1{`RANDOM}};
  FifoCell_244 = _RAND_246[8:0];
  _RAND_247 = {1{`RANDOM}};
  FifoCell_245 = _RAND_247[8:0];
  _RAND_248 = {1{`RANDOM}};
  FifoCell_246 = _RAND_248[8:0];
  _RAND_249 = {1{`RANDOM}};
  FifoCell_247 = _RAND_249[8:0];
  _RAND_250 = {1{`RANDOM}};
  FifoCell_248 = _RAND_250[8:0];
  _RAND_251 = {1{`RANDOM}};
  FifoCell_249 = _RAND_251[8:0];
  _RAND_252 = {1{`RANDOM}};
  FifoCell_250 = _RAND_252[8:0];
  _RAND_253 = {1{`RANDOM}};
  FifoCell_251 = _RAND_253[8:0];
  _RAND_254 = {1{`RANDOM}};
  FifoCell_252 = _RAND_254[8:0];
  _RAND_255 = {1{`RANDOM}};
  FifoCell_253 = _RAND_255[8:0];
  _RAND_256 = {1{`RANDOM}};
  FifoCell_254 = _RAND_256[8:0];
  _RAND_257 = {1{`RANDOM}};
  FifoCell_255 = _RAND_257[8:0];
  _RAND_258 = {1{`RANDOM}};
  FifoCell_256 = _RAND_258[8:0];
  _RAND_259 = {1{`RANDOM}};
  FifoCell_257 = _RAND_259[8:0];
  _RAND_260 = {1{`RANDOM}};
  FifoCell_258 = _RAND_260[8:0];
  _RAND_261 = {1{`RANDOM}};
  FifoCell_259 = _RAND_261[8:0];
  _RAND_262 = {1{`RANDOM}};
  FifoCell_260 = _RAND_262[8:0];
  _RAND_263 = {1{`RANDOM}};
  FifoCell_261 = _RAND_263[8:0];
  _RAND_264 = {1{`RANDOM}};
  FifoCell_262 = _RAND_264[8:0];
  _RAND_265 = {1{`RANDOM}};
  FifoCell_263 = _RAND_265[8:0];
  _RAND_266 = {1{`RANDOM}};
  FifoCell_264 = _RAND_266[8:0];
  _RAND_267 = {1{`RANDOM}};
  FifoCell_265 = _RAND_267[8:0];
  _RAND_268 = {1{`RANDOM}};
  FifoCell_266 = _RAND_268[8:0];
  _RAND_269 = {1{`RANDOM}};
  FifoCell_267 = _RAND_269[8:0];
  _RAND_270 = {1{`RANDOM}};
  FifoCell_268 = _RAND_270[8:0];
  _RAND_271 = {1{`RANDOM}};
  FifoCell_269 = _RAND_271[8:0];
  _RAND_272 = {1{`RANDOM}};
  FifoCell_270 = _RAND_272[8:0];
  _RAND_273 = {1{`RANDOM}};
  FifoCell_271 = _RAND_273[8:0];
  _RAND_274 = {1{`RANDOM}};
  FifoCell_272 = _RAND_274[8:0];
  _RAND_275 = {1{`RANDOM}};
  FifoCell_273 = _RAND_275[8:0];
  _RAND_276 = {1{`RANDOM}};
  FifoCell_274 = _RAND_276[8:0];
  _RAND_277 = {1{`RANDOM}};
  FifoCell_275 = _RAND_277[8:0];
  _RAND_278 = {1{`RANDOM}};
  FifoCell_276 = _RAND_278[8:0];
  _RAND_279 = {1{`RANDOM}};
  FifoCell_277 = _RAND_279[8:0];
  _RAND_280 = {1{`RANDOM}};
  FifoCell_278 = _RAND_280[8:0];
  _RAND_281 = {1{`RANDOM}};
  FifoCell_279 = _RAND_281[8:0];
  _RAND_282 = {1{`RANDOM}};
  FifoCell_280 = _RAND_282[8:0];
  _RAND_283 = {1{`RANDOM}};
  FifoCell_281 = _RAND_283[8:0];
  _RAND_284 = {1{`RANDOM}};
  FifoCell_282 = _RAND_284[8:0];
  _RAND_285 = {1{`RANDOM}};
  FifoCell_283 = _RAND_285[8:0];
  _RAND_286 = {1{`RANDOM}};
  FifoCell_284 = _RAND_286[8:0];
  _RAND_287 = {1{`RANDOM}};
  FifoCell_285 = _RAND_287[8:0];
  _RAND_288 = {1{`RANDOM}};
  FifoCell_286 = _RAND_288[8:0];
  _RAND_289 = {1{`RANDOM}};
  FifoCell_287 = _RAND_289[8:0];
  _RAND_290 = {1{`RANDOM}};
  FifoCell_288 = _RAND_290[8:0];
  _RAND_291 = {1{`RANDOM}};
  FifoCell_289 = _RAND_291[8:0];
  _RAND_292 = {1{`RANDOM}};
  FifoCell_290 = _RAND_292[8:0];
  _RAND_293 = {1{`RANDOM}};
  FifoCell_291 = _RAND_293[8:0];
  _RAND_294 = {1{`RANDOM}};
  FifoCell_292 = _RAND_294[8:0];
  _RAND_295 = {1{`RANDOM}};
  FifoCell_293 = _RAND_295[8:0];
  _RAND_296 = {1{`RANDOM}};
  FifoCell_294 = _RAND_296[8:0];
  _RAND_297 = {1{`RANDOM}};
  FifoCell_295 = _RAND_297[8:0];
  _RAND_298 = {1{`RANDOM}};
  FifoCell_296 = _RAND_298[8:0];
  _RAND_299 = {1{`RANDOM}};
  FifoCell_297 = _RAND_299[8:0];
  _RAND_300 = {1{`RANDOM}};
  FifoCell_298 = _RAND_300[8:0];
  _RAND_301 = {1{`RANDOM}};
  FifoCell_299 = _RAND_301[8:0];
  _RAND_302 = {1{`RANDOM}};
  FifoCell_300 = _RAND_302[8:0];
  _RAND_303 = {1{`RANDOM}};
  FifoCell_301 = _RAND_303[8:0];
  _RAND_304 = {1{`RANDOM}};
  FifoCell_302 = _RAND_304[8:0];
  _RAND_305 = {1{`RANDOM}};
  FifoCell_303 = _RAND_305[8:0];
  _RAND_306 = {1{`RANDOM}};
  FifoCell_304 = _RAND_306[8:0];
  _RAND_307 = {1{`RANDOM}};
  FifoCell_305 = _RAND_307[8:0];
  _RAND_308 = {1{`RANDOM}};
  FifoCell_306 = _RAND_308[8:0];
  _RAND_309 = {1{`RANDOM}};
  FifoCell_307 = _RAND_309[8:0];
  _RAND_310 = {1{`RANDOM}};
  FifoCell_308 = _RAND_310[8:0];
  _RAND_311 = {1{`RANDOM}};
  FifoCell_309 = _RAND_311[8:0];
  _RAND_312 = {1{`RANDOM}};
  FifoCell_310 = _RAND_312[8:0];
  _RAND_313 = {1{`RANDOM}};
  FifoCell_311 = _RAND_313[8:0];
  _RAND_314 = {1{`RANDOM}};
  FifoCell_312 = _RAND_314[8:0];
  _RAND_315 = {1{`RANDOM}};
  FifoCell_313 = _RAND_315[8:0];
  _RAND_316 = {1{`RANDOM}};
  FifoCell_314 = _RAND_316[8:0];
  _RAND_317 = {1{`RANDOM}};
  FifoCell_315 = _RAND_317[8:0];
  _RAND_318 = {1{`RANDOM}};
  FifoCell_316 = _RAND_318[8:0];
  _RAND_319 = {1{`RANDOM}};
  FifoCell_317 = _RAND_319[8:0];
  _RAND_320 = {1{`RANDOM}};
  FifoCell_318 = _RAND_320[8:0];
  _RAND_321 = {1{`RANDOM}};
  FifoCell_319 = _RAND_321[8:0];
  _RAND_322 = {1{`RANDOM}};
  FifoCell_320 = _RAND_322[8:0];
  _RAND_323 = {1{`RANDOM}};
  FifoCell_321 = _RAND_323[8:0];
  _RAND_324 = {1{`RANDOM}};
  FifoCell_322 = _RAND_324[8:0];
  _RAND_325 = {1{`RANDOM}};
  FifoCell_323 = _RAND_325[8:0];
  _RAND_326 = {1{`RANDOM}};
  FifoCell_324 = _RAND_326[8:0];
  _RAND_327 = {1{`RANDOM}};
  FifoCell_325 = _RAND_327[8:0];
  _RAND_328 = {1{`RANDOM}};
  FifoCell_326 = _RAND_328[8:0];
  _RAND_329 = {1{`RANDOM}};
  FifoCell_327 = _RAND_329[8:0];
  _RAND_330 = {1{`RANDOM}};
  FifoCell_328 = _RAND_330[8:0];
  _RAND_331 = {1{`RANDOM}};
  FifoCell_329 = _RAND_331[8:0];
  _RAND_332 = {1{`RANDOM}};
  FifoCell_330 = _RAND_332[8:0];
  _RAND_333 = {1{`RANDOM}};
  FifoCell_331 = _RAND_333[8:0];
  _RAND_334 = {1{`RANDOM}};
  FifoCell_332 = _RAND_334[8:0];
  _RAND_335 = {1{`RANDOM}};
  FifoCell_333 = _RAND_335[8:0];
  _RAND_336 = {1{`RANDOM}};
  FifoCell_334 = _RAND_336[8:0];
  _RAND_337 = {1{`RANDOM}};
  FifoCell_335 = _RAND_337[8:0];
  _RAND_338 = {1{`RANDOM}};
  FifoCell_336 = _RAND_338[8:0];
  _RAND_339 = {1{`RANDOM}};
  FifoCell_337 = _RAND_339[8:0];
  _RAND_340 = {1{`RANDOM}};
  FifoCell_338 = _RAND_340[8:0];
  _RAND_341 = {1{`RANDOM}};
  FifoCell_339 = _RAND_341[8:0];
  _RAND_342 = {1{`RANDOM}};
  FifoCell_340 = _RAND_342[8:0];
  _RAND_343 = {1{`RANDOM}};
  FifoCell_341 = _RAND_343[8:0];
  _RAND_344 = {1{`RANDOM}};
  FifoCell_342 = _RAND_344[8:0];
  _RAND_345 = {1{`RANDOM}};
  FifoCell_343 = _RAND_345[8:0];
  _RAND_346 = {1{`RANDOM}};
  FifoCell_344 = _RAND_346[8:0];
  _RAND_347 = {1{`RANDOM}};
  FifoCell_345 = _RAND_347[8:0];
  _RAND_348 = {1{`RANDOM}};
  FifoCell_346 = _RAND_348[8:0];
  _RAND_349 = {1{`RANDOM}};
  FifoCell_347 = _RAND_349[8:0];
  _RAND_350 = {1{`RANDOM}};
  FifoCell_348 = _RAND_350[8:0];
  _RAND_351 = {1{`RANDOM}};
  FifoCell_349 = _RAND_351[8:0];
  _RAND_352 = {1{`RANDOM}};
  FifoCell_350 = _RAND_352[8:0];
  _RAND_353 = {1{`RANDOM}};
  FifoCell_351 = _RAND_353[8:0];
  _RAND_354 = {1{`RANDOM}};
  FifoCell_352 = _RAND_354[8:0];
  _RAND_355 = {1{`RANDOM}};
  FifoCell_353 = _RAND_355[8:0];
  _RAND_356 = {1{`RANDOM}};
  FifoCell_354 = _RAND_356[8:0];
  _RAND_357 = {1{`RANDOM}};
  FifoCell_355 = _RAND_357[8:0];
  _RAND_358 = {1{`RANDOM}};
  FifoCell_356 = _RAND_358[8:0];
  _RAND_359 = {1{`RANDOM}};
  FifoCell_357 = _RAND_359[8:0];
  _RAND_360 = {1{`RANDOM}};
  FifoCell_358 = _RAND_360[8:0];
  _RAND_361 = {1{`RANDOM}};
  FifoCell_359 = _RAND_361[8:0];
  _RAND_362 = {1{`RANDOM}};
  FifoCell_360 = _RAND_362[8:0];
  _RAND_363 = {1{`RANDOM}};
  FifoCell_361 = _RAND_363[8:0];
  _RAND_364 = {1{`RANDOM}};
  FifoCell_362 = _RAND_364[8:0];
  _RAND_365 = {1{`RANDOM}};
  FifoCell_363 = _RAND_365[8:0];
  _RAND_366 = {1{`RANDOM}};
  FifoCell_364 = _RAND_366[8:0];
  _RAND_367 = {1{`RANDOM}};
  FifoCell_365 = _RAND_367[8:0];
  _RAND_368 = {1{`RANDOM}};
  FifoCell_366 = _RAND_368[8:0];
  _RAND_369 = {1{`RANDOM}};
  FifoCell_367 = _RAND_369[8:0];
  _RAND_370 = {1{`RANDOM}};
  FifoCell_368 = _RAND_370[8:0];
  _RAND_371 = {1{`RANDOM}};
  FifoCell_369 = _RAND_371[8:0];
  _RAND_372 = {1{`RANDOM}};
  FifoCell_370 = _RAND_372[8:0];
  _RAND_373 = {1{`RANDOM}};
  FifoCell_371 = _RAND_373[8:0];
  _RAND_374 = {1{`RANDOM}};
  FifoCell_372 = _RAND_374[8:0];
  _RAND_375 = {1{`RANDOM}};
  FifoCell_373 = _RAND_375[8:0];
  _RAND_376 = {1{`RANDOM}};
  FifoCell_374 = _RAND_376[8:0];
  _RAND_377 = {1{`RANDOM}};
  FifoCell_375 = _RAND_377[8:0];
  _RAND_378 = {1{`RANDOM}};
  FifoCell_376 = _RAND_378[8:0];
  _RAND_379 = {1{`RANDOM}};
  FifoCell_377 = _RAND_379[8:0];
  _RAND_380 = {1{`RANDOM}};
  FifoCell_378 = _RAND_380[8:0];
  _RAND_381 = {1{`RANDOM}};
  FifoCell_379 = _RAND_381[8:0];
  _RAND_382 = {1{`RANDOM}};
  FifoCell_380 = _RAND_382[8:0];
  _RAND_383 = {1{`RANDOM}};
  FifoCell_381 = _RAND_383[8:0];
  _RAND_384 = {1{`RANDOM}};
  FifoCell_382 = _RAND_384[8:0];
  _RAND_385 = {1{`RANDOM}};
  FifoCell_383 = _RAND_385[8:0];
  _RAND_386 = {1{`RANDOM}};
  FifoCell_384 = _RAND_386[8:0];
  _RAND_387 = {1{`RANDOM}};
  FifoCell_385 = _RAND_387[8:0];
  _RAND_388 = {1{`RANDOM}};
  FifoCell_386 = _RAND_388[8:0];
  _RAND_389 = {1{`RANDOM}};
  FifoCell_387 = _RAND_389[8:0];
  _RAND_390 = {1{`RANDOM}};
  FifoCell_388 = _RAND_390[8:0];
  _RAND_391 = {1{`RANDOM}};
  FifoCell_389 = _RAND_391[8:0];
  _RAND_392 = {1{`RANDOM}};
  FifoCell_390 = _RAND_392[8:0];
  _RAND_393 = {1{`RANDOM}};
  FifoCell_391 = _RAND_393[8:0];
  _RAND_394 = {1{`RANDOM}};
  FifoCell_392 = _RAND_394[8:0];
  _RAND_395 = {1{`RANDOM}};
  FifoCell_393 = _RAND_395[8:0];
  _RAND_396 = {1{`RANDOM}};
  FifoCell_394 = _RAND_396[8:0];
  _RAND_397 = {1{`RANDOM}};
  FifoCell_395 = _RAND_397[8:0];
  _RAND_398 = {1{`RANDOM}};
  FifoCell_396 = _RAND_398[8:0];
  _RAND_399 = {1{`RANDOM}};
  FifoCell_397 = _RAND_399[8:0];
  _RAND_400 = {1{`RANDOM}};
  FifoCell_398 = _RAND_400[8:0];
  _RAND_401 = {1{`RANDOM}};
  FifoCell_399 = _RAND_401[8:0];
  _RAND_402 = {1{`RANDOM}};
  FifoCell_400 = _RAND_402[8:0];
  _RAND_403 = {1{`RANDOM}};
  FifoCell_401 = _RAND_403[8:0];
  _RAND_404 = {1{`RANDOM}};
  FifoCell_402 = _RAND_404[8:0];
  _RAND_405 = {1{`RANDOM}};
  FifoCell_403 = _RAND_405[8:0];
  _RAND_406 = {1{`RANDOM}};
  FifoCell_404 = _RAND_406[8:0];
  _RAND_407 = {1{`RANDOM}};
  FifoCell_405 = _RAND_407[8:0];
  _RAND_408 = {1{`RANDOM}};
  FifoCell_406 = _RAND_408[8:0];
  _RAND_409 = {1{`RANDOM}};
  FifoCell_407 = _RAND_409[8:0];
  _RAND_410 = {1{`RANDOM}};
  FifoCell_408 = _RAND_410[8:0];
  _RAND_411 = {1{`RANDOM}};
  FifoCell_409 = _RAND_411[8:0];
  _RAND_412 = {1{`RANDOM}};
  FifoCell_410 = _RAND_412[8:0];
  _RAND_413 = {1{`RANDOM}};
  FifoCell_411 = _RAND_413[8:0];
  _RAND_414 = {1{`RANDOM}};
  FifoCell_412 = _RAND_414[8:0];
  _RAND_415 = {1{`RANDOM}};
  FifoCell_413 = _RAND_415[8:0];
  _RAND_416 = {1{`RANDOM}};
  FifoCell_414 = _RAND_416[8:0];
  _RAND_417 = {1{`RANDOM}};
  FifoCell_415 = _RAND_417[8:0];
  _RAND_418 = {1{`RANDOM}};
  FifoCell_416 = _RAND_418[8:0];
  _RAND_419 = {1{`RANDOM}};
  FifoCell_417 = _RAND_419[8:0];
  _RAND_420 = {1{`RANDOM}};
  FifoCell_418 = _RAND_420[8:0];
  _RAND_421 = {1{`RANDOM}};
  FifoCell_419 = _RAND_421[8:0];
  _RAND_422 = {1{`RANDOM}};
  FifoCell_420 = _RAND_422[8:0];
  _RAND_423 = {1{`RANDOM}};
  FifoCell_421 = _RAND_423[8:0];
  _RAND_424 = {1{`RANDOM}};
  FifoCell_422 = _RAND_424[8:0];
  _RAND_425 = {1{`RANDOM}};
  FifoCell_423 = _RAND_425[8:0];
  _RAND_426 = {1{`RANDOM}};
  FifoCell_424 = _RAND_426[8:0];
  _RAND_427 = {1{`RANDOM}};
  FifoCell_425 = _RAND_427[8:0];
  _RAND_428 = {1{`RANDOM}};
  FifoCell_426 = _RAND_428[8:0];
  _RAND_429 = {1{`RANDOM}};
  FifoCell_427 = _RAND_429[8:0];
  _RAND_430 = {1{`RANDOM}};
  FifoCell_428 = _RAND_430[8:0];
  _RAND_431 = {1{`RANDOM}};
  FifoCell_429 = _RAND_431[8:0];
  _RAND_432 = {1{`RANDOM}};
  FifoCell_430 = _RAND_432[8:0];
  _RAND_433 = {1{`RANDOM}};
  FifoCell_431 = _RAND_433[8:0];
  _RAND_434 = {1{`RANDOM}};
  FifoCell_432 = _RAND_434[8:0];
  _RAND_435 = {1{`RANDOM}};
  FifoCell_433 = _RAND_435[8:0];
  _RAND_436 = {1{`RANDOM}};
  FifoCell_434 = _RAND_436[8:0];
  _RAND_437 = {1{`RANDOM}};
  FifoCell_435 = _RAND_437[8:0];
  _RAND_438 = {1{`RANDOM}};
  FifoCell_436 = _RAND_438[8:0];
  _RAND_439 = {1{`RANDOM}};
  FifoCell_437 = _RAND_439[8:0];
  _RAND_440 = {1{`RANDOM}};
  FifoCell_438 = _RAND_440[8:0];
  _RAND_441 = {1{`RANDOM}};
  FifoCell_439 = _RAND_441[8:0];
  _RAND_442 = {1{`RANDOM}};
  FifoCell_440 = _RAND_442[8:0];
  _RAND_443 = {1{`RANDOM}};
  FifoCell_441 = _RAND_443[8:0];
  _RAND_444 = {1{`RANDOM}};
  FifoCell_442 = _RAND_444[8:0];
  _RAND_445 = {1{`RANDOM}};
  FifoCell_443 = _RAND_445[8:0];
  _RAND_446 = {1{`RANDOM}};
  FifoCell_444 = _RAND_446[8:0];
  _RAND_447 = {1{`RANDOM}};
  FifoCell_445 = _RAND_447[8:0];
  _RAND_448 = {1{`RANDOM}};
  FifoCell_446 = _RAND_448[8:0];
  _RAND_449 = {1{`RANDOM}};
  FifoCell_447 = _RAND_449[8:0];
  _RAND_450 = {1{`RANDOM}};
  FifoCell_448 = _RAND_450[8:0];
  _RAND_451 = {1{`RANDOM}};
  FifoCell_449 = _RAND_451[8:0];
  _RAND_452 = {1{`RANDOM}};
  FifoCell_450 = _RAND_452[8:0];
  _RAND_453 = {1{`RANDOM}};
  FifoCell_451 = _RAND_453[8:0];
  _RAND_454 = {1{`RANDOM}};
  FifoCell_452 = _RAND_454[8:0];
  _RAND_455 = {1{`RANDOM}};
  FifoCell_453 = _RAND_455[8:0];
  _RAND_456 = {1{`RANDOM}};
  FifoCell_454 = _RAND_456[8:0];
  _RAND_457 = {1{`RANDOM}};
  FifoCell_455 = _RAND_457[8:0];
  _RAND_458 = {1{`RANDOM}};
  FifoCell_456 = _RAND_458[8:0];
  _RAND_459 = {1{`RANDOM}};
  FifoCell_457 = _RAND_459[8:0];
  _RAND_460 = {1{`RANDOM}};
  FifoCell_458 = _RAND_460[8:0];
  _RAND_461 = {1{`RANDOM}};
  FifoCell_459 = _RAND_461[8:0];
  _RAND_462 = {1{`RANDOM}};
  FifoCell_460 = _RAND_462[8:0];
  _RAND_463 = {1{`RANDOM}};
  FifoCell_461 = _RAND_463[8:0];
  _RAND_464 = {1{`RANDOM}};
  FifoCell_462 = _RAND_464[8:0];
  _RAND_465 = {1{`RANDOM}};
  FifoCell_463 = _RAND_465[8:0];
  _RAND_466 = {1{`RANDOM}};
  FifoCell_464 = _RAND_466[8:0];
  _RAND_467 = {1{`RANDOM}};
  FifoCell_465 = _RAND_467[8:0];
  _RAND_468 = {1{`RANDOM}};
  FifoCell_466 = _RAND_468[8:0];
  _RAND_469 = {1{`RANDOM}};
  FifoCell_467 = _RAND_469[8:0];
  _RAND_470 = {1{`RANDOM}};
  FifoCell_468 = _RAND_470[8:0];
  _RAND_471 = {1{`RANDOM}};
  FifoCell_469 = _RAND_471[8:0];
  _RAND_472 = {1{`RANDOM}};
  FifoCell_470 = _RAND_472[8:0];
  _RAND_473 = {1{`RANDOM}};
  FifoCell_471 = _RAND_473[8:0];
  _RAND_474 = {1{`RANDOM}};
  FifoCell_472 = _RAND_474[8:0];
  _RAND_475 = {1{`RANDOM}};
  FifoCell_473 = _RAND_475[8:0];
  _RAND_476 = {1{`RANDOM}};
  FifoCell_474 = _RAND_476[8:0];
  _RAND_477 = {1{`RANDOM}};
  FifoCell_475 = _RAND_477[8:0];
  _RAND_478 = {1{`RANDOM}};
  FifoCell_476 = _RAND_478[8:0];
  _RAND_479 = {1{`RANDOM}};
  FifoCell_477 = _RAND_479[8:0];
  _RAND_480 = {1{`RANDOM}};
  FifoCell_478 = _RAND_480[8:0];
  _RAND_481 = {1{`RANDOM}};
  FifoCell_479 = _RAND_481[8:0];
  _RAND_482 = {1{`RANDOM}};
  FifoCell_480 = _RAND_482[8:0];
  _RAND_483 = {1{`RANDOM}};
  FifoCell_481 = _RAND_483[8:0];
  _RAND_484 = {1{`RANDOM}};
  FifoCell_482 = _RAND_484[8:0];
  _RAND_485 = {1{`RANDOM}};
  FifoCell_483 = _RAND_485[8:0];
  _RAND_486 = {1{`RANDOM}};
  FifoCell_484 = _RAND_486[8:0];
  _RAND_487 = {1{`RANDOM}};
  FifoCell_485 = _RAND_487[8:0];
  _RAND_488 = {1{`RANDOM}};
  FifoCell_486 = _RAND_488[8:0];
  _RAND_489 = {1{`RANDOM}};
  FifoCell_487 = _RAND_489[8:0];
  _RAND_490 = {1{`RANDOM}};
  FifoCell_488 = _RAND_490[8:0];
  _RAND_491 = {1{`RANDOM}};
  FifoCell_489 = _RAND_491[8:0];
  _RAND_492 = {1{`RANDOM}};
  FifoCell_490 = _RAND_492[8:0];
  _RAND_493 = {1{`RANDOM}};
  FifoCell_491 = _RAND_493[8:0];
  _RAND_494 = {1{`RANDOM}};
  FifoCell_492 = _RAND_494[8:0];
  _RAND_495 = {1{`RANDOM}};
  FifoCell_493 = _RAND_495[8:0];
  _RAND_496 = {1{`RANDOM}};
  FifoCell_494 = _RAND_496[8:0];
  _RAND_497 = {1{`RANDOM}};
  FifoCell_495 = _RAND_497[8:0];
  _RAND_498 = {1{`RANDOM}};
  FifoCell_496 = _RAND_498[8:0];
  _RAND_499 = {1{`RANDOM}};
  FifoCell_497 = _RAND_499[8:0];
  _RAND_500 = {1{`RANDOM}};
  FifoCell_498 = _RAND_500[8:0];
  _RAND_501 = {1{`RANDOM}};
  FifoCell_499 = _RAND_501[8:0];
  _RAND_502 = {1{`RANDOM}};
  FifoCell_500 = _RAND_502[8:0];
  _RAND_503 = {1{`RANDOM}};
  FifoCell_501 = _RAND_503[8:0];
  _RAND_504 = {1{`RANDOM}};
  FifoCell_502 = _RAND_504[8:0];
  _RAND_505 = {1{`RANDOM}};
  FifoCell_503 = _RAND_505[8:0];
  _RAND_506 = {1{`RANDOM}};
  FifoCell_504 = _RAND_506[8:0];
  _RAND_507 = {1{`RANDOM}};
  FifoCell_505 = _RAND_507[8:0];
  _RAND_508 = {1{`RANDOM}};
  FifoCell_506 = _RAND_508[8:0];
  _RAND_509 = {1{`RANDOM}};
  FifoCell_507 = _RAND_509[8:0];
  _RAND_510 = {1{`RANDOM}};
  FifoCell_508 = _RAND_510[8:0];
  _RAND_511 = {1{`RANDOM}};
  FifoCell_509 = _RAND_511[8:0];
  _RAND_512 = {1{`RANDOM}};
  FifoCell_510 = _RAND_512[8:0];
  _RAND_513 = {1{`RANDOM}};
  FifoCell_511 = _RAND_513[8:0];
  _RAND_514 = {1{`RANDOM}};
  FifoCell_512 = _RAND_514[8:0];
  _RAND_515 = {1{`RANDOM}};
  FifoCell_513 = _RAND_515[8:0];
  _RAND_516 = {1{`RANDOM}};
  FifoCell_514 = _RAND_516[8:0];
  _RAND_517 = {1{`RANDOM}};
  FifoCell_515 = _RAND_517[8:0];
  _RAND_518 = {1{`RANDOM}};
  FifoCell_516 = _RAND_518[8:0];
  _RAND_519 = {1{`RANDOM}};
  FifoCell_517 = _RAND_519[8:0];
  _RAND_520 = {1{`RANDOM}};
  FifoCell_518 = _RAND_520[8:0];
  _RAND_521 = {1{`RANDOM}};
  FifoCell_519 = _RAND_521[8:0];
  _RAND_522 = {1{`RANDOM}};
  FifoCell_520 = _RAND_522[8:0];
  _RAND_523 = {1{`RANDOM}};
  FifoCell_521 = _RAND_523[8:0];
  _RAND_524 = {1{`RANDOM}};
  FifoCell_522 = _RAND_524[8:0];
  _RAND_525 = {1{`RANDOM}};
  FifoCell_523 = _RAND_525[8:0];
  _RAND_526 = {1{`RANDOM}};
  FifoCell_524 = _RAND_526[8:0];
  _RAND_527 = {1{`RANDOM}};
  FifoCell_525 = _RAND_527[8:0];
  _RAND_528 = {1{`RANDOM}};
  FifoCell_526 = _RAND_528[8:0];
  _RAND_529 = {1{`RANDOM}};
  FifoCell_527 = _RAND_529[8:0];
  _RAND_530 = {1{`RANDOM}};
  FifoCell_528 = _RAND_530[8:0];
  _RAND_531 = {1{`RANDOM}};
  FifoCell_529 = _RAND_531[8:0];
  _RAND_532 = {1{`RANDOM}};
  FifoCell_530 = _RAND_532[8:0];
  _RAND_533 = {1{`RANDOM}};
  FifoCell_531 = _RAND_533[8:0];
  _RAND_534 = {1{`RANDOM}};
  FifoCell_532 = _RAND_534[8:0];
  _RAND_535 = {1{`RANDOM}};
  FifoCell_533 = _RAND_535[8:0];
  _RAND_536 = {1{`RANDOM}};
  FifoCell_534 = _RAND_536[8:0];
  _RAND_537 = {1{`RANDOM}};
  FifoCell_535 = _RAND_537[8:0];
  _RAND_538 = {1{`RANDOM}};
  FifoCell_536 = _RAND_538[8:0];
  _RAND_539 = {1{`RANDOM}};
  FifoCell_537 = _RAND_539[8:0];
  _RAND_540 = {1{`RANDOM}};
  FifoCell_538 = _RAND_540[8:0];
  _RAND_541 = {1{`RANDOM}};
  FifoCell_539 = _RAND_541[8:0];
  _RAND_542 = {1{`RANDOM}};
  FifoCell_540 = _RAND_542[8:0];
  _RAND_543 = {1{`RANDOM}};
  FifoCell_541 = _RAND_543[8:0];
  _RAND_544 = {1{`RANDOM}};
  FifoCell_542 = _RAND_544[8:0];
  _RAND_545 = {1{`RANDOM}};
  FifoCell_543 = _RAND_545[8:0];
  _RAND_546 = {1{`RANDOM}};
  FifoCell_544 = _RAND_546[8:0];
  _RAND_547 = {1{`RANDOM}};
  FifoCell_545 = _RAND_547[8:0];
  _RAND_548 = {1{`RANDOM}};
  FifoCell_546 = _RAND_548[8:0];
  _RAND_549 = {1{`RANDOM}};
  FifoCell_547 = _RAND_549[8:0];
  _RAND_550 = {1{`RANDOM}};
  FifoCell_548 = _RAND_550[8:0];
  _RAND_551 = {1{`RANDOM}};
  FifoCell_549 = _RAND_551[8:0];
  _RAND_552 = {1{`RANDOM}};
  FifoCell_550 = _RAND_552[8:0];
  _RAND_553 = {1{`RANDOM}};
  FifoCell_551 = _RAND_553[8:0];
  _RAND_554 = {1{`RANDOM}};
  FifoCell_552 = _RAND_554[8:0];
  _RAND_555 = {1{`RANDOM}};
  FifoCell_553 = _RAND_555[8:0];
  _RAND_556 = {1{`RANDOM}};
  FifoCell_554 = _RAND_556[8:0];
  _RAND_557 = {1{`RANDOM}};
  FifoCell_555 = _RAND_557[8:0];
  _RAND_558 = {1{`RANDOM}};
  FifoCell_556 = _RAND_558[8:0];
  _RAND_559 = {1{`RANDOM}};
  FifoCell_557 = _RAND_559[8:0];
  _RAND_560 = {1{`RANDOM}};
  FifoCell_558 = _RAND_560[8:0];
  _RAND_561 = {1{`RANDOM}};
  FifoCell_559 = _RAND_561[8:0];
  _RAND_562 = {1{`RANDOM}};
  FifoCell_560 = _RAND_562[8:0];
  _RAND_563 = {1{`RANDOM}};
  FifoCell_561 = _RAND_563[8:0];
  _RAND_564 = {1{`RANDOM}};
  FifoCell_562 = _RAND_564[8:0];
  _RAND_565 = {1{`RANDOM}};
  FifoCell_563 = _RAND_565[8:0];
  _RAND_566 = {1{`RANDOM}};
  FifoCell_564 = _RAND_566[8:0];
  _RAND_567 = {1{`RANDOM}};
  FifoCell_565 = _RAND_567[8:0];
  _RAND_568 = {1{`RANDOM}};
  FifoCell_566 = _RAND_568[8:0];
  _RAND_569 = {1{`RANDOM}};
  FifoCell_567 = _RAND_569[8:0];
  _RAND_570 = {1{`RANDOM}};
  FifoCell_568 = _RAND_570[8:0];
  _RAND_571 = {1{`RANDOM}};
  FifoCell_569 = _RAND_571[8:0];
  _RAND_572 = {1{`RANDOM}};
  FifoCell_570 = _RAND_572[8:0];
  _RAND_573 = {1{`RANDOM}};
  FifoCell_571 = _RAND_573[8:0];
  _RAND_574 = {1{`RANDOM}};
  FifoCell_572 = _RAND_574[8:0];
  _RAND_575 = {1{`RANDOM}};
  FifoCell_573 = _RAND_575[8:0];
  _RAND_576 = {1{`RANDOM}};
  FifoCell_574 = _RAND_576[8:0];
  _RAND_577 = {1{`RANDOM}};
  FifoCell_575 = _RAND_577[8:0];
  _RAND_578 = {1{`RANDOM}};
  FifoCell_576 = _RAND_578[8:0];
  _RAND_579 = {1{`RANDOM}};
  FifoCell_577 = _RAND_579[8:0];
  _RAND_580 = {1{`RANDOM}};
  FifoCell_578 = _RAND_580[8:0];
  _RAND_581 = {1{`RANDOM}};
  FifoCell_579 = _RAND_581[8:0];
  _RAND_582 = {1{`RANDOM}};
  FifoCell_580 = _RAND_582[8:0];
  _RAND_583 = {1{`RANDOM}};
  FifoCell_581 = _RAND_583[8:0];
  _RAND_584 = {1{`RANDOM}};
  FifoCell_582 = _RAND_584[8:0];
  _RAND_585 = {1{`RANDOM}};
  FifoCell_583 = _RAND_585[8:0];
  _RAND_586 = {1{`RANDOM}};
  FifoCell_584 = _RAND_586[8:0];
  _RAND_587 = {1{`RANDOM}};
  FifoCell_585 = _RAND_587[8:0];
  _RAND_588 = {1{`RANDOM}};
  FifoCell_586 = _RAND_588[8:0];
  _RAND_589 = {1{`RANDOM}};
  FifoCell_587 = _RAND_589[8:0];
  _RAND_590 = {1{`RANDOM}};
  FifoCell_588 = _RAND_590[8:0];
  _RAND_591 = {1{`RANDOM}};
  FifoCell_589 = _RAND_591[8:0];
  _RAND_592 = {1{`RANDOM}};
  FifoCell_590 = _RAND_592[8:0];
  _RAND_593 = {1{`RANDOM}};
  FifoCell_591 = _RAND_593[8:0];
  _RAND_594 = {1{`RANDOM}};
  FifoCell_592 = _RAND_594[8:0];
  _RAND_595 = {1{`RANDOM}};
  FifoCell_593 = _RAND_595[8:0];
  _RAND_596 = {1{`RANDOM}};
  FifoCell_594 = _RAND_596[8:0];
  _RAND_597 = {1{`RANDOM}};
  FifoCell_595 = _RAND_597[8:0];
  _RAND_598 = {1{`RANDOM}};
  FifoCell_596 = _RAND_598[8:0];
  _RAND_599 = {1{`RANDOM}};
  FifoCell_597 = _RAND_599[8:0];
  _RAND_600 = {1{`RANDOM}};
  FifoCell_598 = _RAND_600[8:0];
  _RAND_601 = {1{`RANDOM}};
  FifoCell_599 = _RAND_601[8:0];
  _RAND_602 = {1{`RANDOM}};
  FifoCell_600 = _RAND_602[8:0];
  _RAND_603 = {1{`RANDOM}};
  FifoCell_601 = _RAND_603[8:0];
  _RAND_604 = {1{`RANDOM}};
  FifoCell_602 = _RAND_604[8:0];
  _RAND_605 = {1{`RANDOM}};
  FifoCell_603 = _RAND_605[8:0];
  _RAND_606 = {1{`RANDOM}};
  FifoCell_604 = _RAND_606[8:0];
  _RAND_607 = {1{`RANDOM}};
  FifoCell_605 = _RAND_607[8:0];
  _RAND_608 = {1{`RANDOM}};
  FifoCell_606 = _RAND_608[8:0];
  _RAND_609 = {1{`RANDOM}};
  FifoCell_607 = _RAND_609[8:0];
  _RAND_610 = {1{`RANDOM}};
  FifoCell_608 = _RAND_610[8:0];
  _RAND_611 = {1{`RANDOM}};
  FifoCell_609 = _RAND_611[8:0];
  _RAND_612 = {1{`RANDOM}};
  FifoCell_610 = _RAND_612[8:0];
  _RAND_613 = {1{`RANDOM}};
  FifoCell_611 = _RAND_613[8:0];
  _RAND_614 = {1{`RANDOM}};
  FifoCell_612 = _RAND_614[8:0];
  _RAND_615 = {1{`RANDOM}};
  FifoCell_613 = _RAND_615[8:0];
  _RAND_616 = {1{`RANDOM}};
  FifoCell_614 = _RAND_616[8:0];
  _RAND_617 = {1{`RANDOM}};
  FifoCell_615 = _RAND_617[8:0];
  _RAND_618 = {1{`RANDOM}};
  FifoCell_616 = _RAND_618[8:0];
  _RAND_619 = {1{`RANDOM}};
  FifoCell_617 = _RAND_619[8:0];
  _RAND_620 = {1{`RANDOM}};
  FifoCell_618 = _RAND_620[8:0];
  _RAND_621 = {1{`RANDOM}};
  FifoCell_619 = _RAND_621[8:0];
  _RAND_622 = {1{`RANDOM}};
  FifoCell_620 = _RAND_622[8:0];
  _RAND_623 = {1{`RANDOM}};
  FifoCell_621 = _RAND_623[8:0];
  _RAND_624 = {1{`RANDOM}};
  FifoCell_622 = _RAND_624[8:0];
  _RAND_625 = {1{`RANDOM}};
  FifoCell_623 = _RAND_625[8:0];
  _RAND_626 = {1{`RANDOM}};
  FifoCell_624 = _RAND_626[8:0];
  _RAND_627 = {1{`RANDOM}};
  FifoCell_625 = _RAND_627[8:0];
  _RAND_628 = {1{`RANDOM}};
  FifoCell_626 = _RAND_628[8:0];
  _RAND_629 = {1{`RANDOM}};
  FifoCell_627 = _RAND_629[8:0];
  _RAND_630 = {1{`RANDOM}};
  FifoCell_628 = _RAND_630[8:0];
  _RAND_631 = {1{`RANDOM}};
  FifoCell_629 = _RAND_631[8:0];
  _RAND_632 = {1{`RANDOM}};
  FifoCell_630 = _RAND_632[8:0];
  _RAND_633 = {1{`RANDOM}};
  FifoCell_631 = _RAND_633[8:0];
  _RAND_634 = {1{`RANDOM}};
  FifoCell_632 = _RAND_634[8:0];
  _RAND_635 = {1{`RANDOM}};
  FifoCell_633 = _RAND_635[8:0];
  _RAND_636 = {1{`RANDOM}};
  FifoCell_634 = _RAND_636[8:0];
  _RAND_637 = {1{`RANDOM}};
  FifoCell_635 = _RAND_637[8:0];
  _RAND_638 = {1{`RANDOM}};
  FifoCell_636 = _RAND_638[8:0];
  _RAND_639 = {1{`RANDOM}};
  FifoCell_637 = _RAND_639[8:0];
  _RAND_640 = {1{`RANDOM}};
  FifoCell_638 = _RAND_640[8:0];
  _RAND_641 = {1{`RANDOM}};
  FifoCell_639 = _RAND_641[8:0];
  _RAND_642 = {1{`RANDOM}};
  FifoCell_640 = _RAND_642[8:0];
  _RAND_643 = {1{`RANDOM}};
  FifoCell_641 = _RAND_643[8:0];
  _RAND_644 = {1{`RANDOM}};
  FifoCell_642 = _RAND_644[8:0];
  _RAND_645 = {1{`RANDOM}};
  FifoCell_643 = _RAND_645[8:0];
  _RAND_646 = {1{`RANDOM}};
  FifoCell_644 = _RAND_646[8:0];
  _RAND_647 = {1{`RANDOM}};
  FifoCell_645 = _RAND_647[8:0];
  _RAND_648 = {1{`RANDOM}};
  FifoCell_646 = _RAND_648[8:0];
  _RAND_649 = {1{`RANDOM}};
  FifoCell_647 = _RAND_649[8:0];
  _RAND_650 = {1{`RANDOM}};
  FifoCell_648 = _RAND_650[8:0];
  _RAND_651 = {1{`RANDOM}};
  FifoCell_649 = _RAND_651[8:0];
  _RAND_652 = {1{`RANDOM}};
  FifoCell_650 = _RAND_652[8:0];
  _RAND_653 = {1{`RANDOM}};
  FifoCell_651 = _RAND_653[8:0];
  _RAND_654 = {1{`RANDOM}};
  FifoCell_652 = _RAND_654[8:0];
  _RAND_655 = {1{`RANDOM}};
  FifoCell_653 = _RAND_655[8:0];
  _RAND_656 = {1{`RANDOM}};
  FifoCell_654 = _RAND_656[8:0];
  _RAND_657 = {1{`RANDOM}};
  FifoCell_655 = _RAND_657[8:0];
  _RAND_658 = {1{`RANDOM}};
  FifoCell_656 = _RAND_658[8:0];
  _RAND_659 = {1{`RANDOM}};
  FifoCell_657 = _RAND_659[8:0];
  _RAND_660 = {1{`RANDOM}};
  FifoCell_658 = _RAND_660[8:0];
  _RAND_661 = {1{`RANDOM}};
  FifoCell_659 = _RAND_661[8:0];
  _RAND_662 = {1{`RANDOM}};
  FifoCell_660 = _RAND_662[8:0];
  _RAND_663 = {1{`RANDOM}};
  FifoCell_661 = _RAND_663[8:0];
  _RAND_664 = {1{`RANDOM}};
  FifoCell_662 = _RAND_664[8:0];
  _RAND_665 = {1{`RANDOM}};
  FifoCell_663 = _RAND_665[8:0];
  _RAND_666 = {1{`RANDOM}};
  FifoCell_664 = _RAND_666[8:0];
  _RAND_667 = {1{`RANDOM}};
  FifoCell_665 = _RAND_667[8:0];
  _RAND_668 = {1{`RANDOM}};
  FifoCell_666 = _RAND_668[8:0];
  _RAND_669 = {1{`RANDOM}};
  FifoCell_667 = _RAND_669[8:0];
  _RAND_670 = {1{`RANDOM}};
  FifoCell_668 = _RAND_670[8:0];
  _RAND_671 = {1{`RANDOM}};
  FifoCell_669 = _RAND_671[8:0];
  _RAND_672 = {1{`RANDOM}};
  FifoCell_670 = _RAND_672[8:0];
  _RAND_673 = {1{`RANDOM}};
  FifoCell_671 = _RAND_673[8:0];
  _RAND_674 = {1{`RANDOM}};
  FifoCell_672 = _RAND_674[8:0];
  _RAND_675 = {1{`RANDOM}};
  FifoCell_673 = _RAND_675[8:0];
  _RAND_676 = {1{`RANDOM}};
  FifoCell_674 = _RAND_676[8:0];
  _RAND_677 = {1{`RANDOM}};
  FifoCell_675 = _RAND_677[8:0];
  _RAND_678 = {1{`RANDOM}};
  FifoCell_676 = _RAND_678[8:0];
  _RAND_679 = {1{`RANDOM}};
  FifoCell_677 = _RAND_679[8:0];
  _RAND_680 = {1{`RANDOM}};
  FifoCell_678 = _RAND_680[8:0];
  _RAND_681 = {1{`RANDOM}};
  FifoCell_679 = _RAND_681[8:0];
  _RAND_682 = {1{`RANDOM}};
  FifoCell_680 = _RAND_682[8:0];
  _RAND_683 = {1{`RANDOM}};
  FifoCell_681 = _RAND_683[8:0];
  _RAND_684 = {1{`RANDOM}};
  FifoCell_682 = _RAND_684[8:0];
  _RAND_685 = {1{`RANDOM}};
  FifoCell_683 = _RAND_685[8:0];
  _RAND_686 = {1{`RANDOM}};
  FifoCell_684 = _RAND_686[8:0];
  _RAND_687 = {1{`RANDOM}};
  FifoCell_685 = _RAND_687[8:0];
  _RAND_688 = {1{`RANDOM}};
  FifoCell_686 = _RAND_688[8:0];
  _RAND_689 = {1{`RANDOM}};
  FifoCell_687 = _RAND_689[8:0];
  _RAND_690 = {1{`RANDOM}};
  FifoCell_688 = _RAND_690[8:0];
  _RAND_691 = {1{`RANDOM}};
  FifoCell_689 = _RAND_691[8:0];
  _RAND_692 = {1{`RANDOM}};
  FifoCell_690 = _RAND_692[8:0];
  _RAND_693 = {1{`RANDOM}};
  FifoCell_691 = _RAND_693[8:0];
  _RAND_694 = {1{`RANDOM}};
  FifoCell_692 = _RAND_694[8:0];
  _RAND_695 = {1{`RANDOM}};
  FifoCell_693 = _RAND_695[8:0];
  _RAND_696 = {1{`RANDOM}};
  FifoCell_694 = _RAND_696[8:0];
  _RAND_697 = {1{`RANDOM}};
  FifoCell_695 = _RAND_697[8:0];
  _RAND_698 = {1{`RANDOM}};
  FifoCell_696 = _RAND_698[8:0];
  _RAND_699 = {1{`RANDOM}};
  FifoCell_697 = _RAND_699[8:0];
  _RAND_700 = {1{`RANDOM}};
  FifoCell_698 = _RAND_700[8:0];
  _RAND_701 = {1{`RANDOM}};
  FifoCell_699 = _RAND_701[8:0];
  _RAND_702 = {1{`RANDOM}};
  FifoCell_700 = _RAND_702[8:0];
  _RAND_703 = {1{`RANDOM}};
  FifoCell_701 = _RAND_703[8:0];
  _RAND_704 = {1{`RANDOM}};
  FifoCell_702 = _RAND_704[8:0];
  _RAND_705 = {1{`RANDOM}};
  FifoCell_703 = _RAND_705[8:0];
  _RAND_706 = {1{`RANDOM}};
  FifoCell_704 = _RAND_706[8:0];
  _RAND_707 = {1{`RANDOM}};
  FifoCell_705 = _RAND_707[8:0];
  _RAND_708 = {1{`RANDOM}};
  FifoCell_706 = _RAND_708[8:0];
  _RAND_709 = {1{`RANDOM}};
  FifoCell_707 = _RAND_709[8:0];
  _RAND_710 = {1{`RANDOM}};
  FifoCell_708 = _RAND_710[8:0];
  _RAND_711 = {1{`RANDOM}};
  FifoCell_709 = _RAND_711[8:0];
  _RAND_712 = {1{`RANDOM}};
  FifoCell_710 = _RAND_712[8:0];
  _RAND_713 = {1{`RANDOM}};
  FifoCell_711 = _RAND_713[8:0];
  _RAND_714 = {1{`RANDOM}};
  FifoCell_712 = _RAND_714[8:0];
  _RAND_715 = {1{`RANDOM}};
  FifoCell_713 = _RAND_715[8:0];
  _RAND_716 = {1{`RANDOM}};
  FifoCell_714 = _RAND_716[8:0];
  _RAND_717 = {1{`RANDOM}};
  FifoCell_715 = _RAND_717[8:0];
  _RAND_718 = {1{`RANDOM}};
  FifoCell_716 = _RAND_718[8:0];
  _RAND_719 = {1{`RANDOM}};
  FifoCell_717 = _RAND_719[8:0];
  _RAND_720 = {1{`RANDOM}};
  FifoCell_718 = _RAND_720[8:0];
  _RAND_721 = {1{`RANDOM}};
  FifoCell_719 = _RAND_721[8:0];
  _RAND_722 = {1{`RANDOM}};
  FifoCell_720 = _RAND_722[8:0];
  _RAND_723 = {1{`RANDOM}};
  FifoCell_721 = _RAND_723[8:0];
  _RAND_724 = {1{`RANDOM}};
  FifoCell_722 = _RAND_724[8:0];
  _RAND_725 = {1{`RANDOM}};
  FifoCell_723 = _RAND_725[8:0];
  _RAND_726 = {1{`RANDOM}};
  FifoCell_724 = _RAND_726[8:0];
  _RAND_727 = {1{`RANDOM}};
  FifoCell_725 = _RAND_727[8:0];
  _RAND_728 = {1{`RANDOM}};
  FifoCell_726 = _RAND_728[8:0];
  _RAND_729 = {1{`RANDOM}};
  FifoCell_727 = _RAND_729[8:0];
  _RAND_730 = {1{`RANDOM}};
  FifoCell_728 = _RAND_730[8:0];
  _RAND_731 = {1{`RANDOM}};
  FifoCell_729 = _RAND_731[8:0];
  _RAND_732 = {1{`RANDOM}};
  FifoCell_730 = _RAND_732[8:0];
  _RAND_733 = {1{`RANDOM}};
  FifoCell_731 = _RAND_733[8:0];
  _RAND_734 = {1{`RANDOM}};
  FifoCell_732 = _RAND_734[8:0];
  _RAND_735 = {1{`RANDOM}};
  FifoCell_733 = _RAND_735[8:0];
  _RAND_736 = {1{`RANDOM}};
  FifoCell_734 = _RAND_736[8:0];
  _RAND_737 = {1{`RANDOM}};
  FifoCell_735 = _RAND_737[8:0];
  _RAND_738 = {1{`RANDOM}};
  FifoCell_736 = _RAND_738[8:0];
  _RAND_739 = {1{`RANDOM}};
  FifoCell_737 = _RAND_739[8:0];
  _RAND_740 = {1{`RANDOM}};
  FifoCell_738 = _RAND_740[8:0];
  _RAND_741 = {1{`RANDOM}};
  FifoCell_739 = _RAND_741[8:0];
  _RAND_742 = {1{`RANDOM}};
  FifoCell_740 = _RAND_742[8:0];
  _RAND_743 = {1{`RANDOM}};
  FifoCell_741 = _RAND_743[8:0];
  _RAND_744 = {1{`RANDOM}};
  FifoCell_742 = _RAND_744[8:0];
  _RAND_745 = {1{`RANDOM}};
  FifoCell_743 = _RAND_745[8:0];
  _RAND_746 = {1{`RANDOM}};
  FifoCell_744 = _RAND_746[8:0];
  _RAND_747 = {1{`RANDOM}};
  FifoCell_745 = _RAND_747[8:0];
  _RAND_748 = {1{`RANDOM}};
  FifoCell_746 = _RAND_748[8:0];
  _RAND_749 = {1{`RANDOM}};
  FifoCell_747 = _RAND_749[8:0];
  _RAND_750 = {1{`RANDOM}};
  FifoCell_748 = _RAND_750[8:0];
  _RAND_751 = {1{`RANDOM}};
  FifoCell_749 = _RAND_751[8:0];
  _RAND_752 = {1{`RANDOM}};
  FifoCell_750 = _RAND_752[8:0];
  _RAND_753 = {1{`RANDOM}};
  FifoCell_751 = _RAND_753[8:0];
  _RAND_754 = {1{`RANDOM}};
  FifoCell_752 = _RAND_754[8:0];
  _RAND_755 = {1{`RANDOM}};
  FifoCell_753 = _RAND_755[8:0];
  _RAND_756 = {1{`RANDOM}};
  FifoCell_754 = _RAND_756[8:0];
  _RAND_757 = {1{`RANDOM}};
  FifoCell_755 = _RAND_757[8:0];
  _RAND_758 = {1{`RANDOM}};
  FifoCell_756 = _RAND_758[8:0];
  _RAND_759 = {1{`RANDOM}};
  FifoCell_757 = _RAND_759[8:0];
  _RAND_760 = {1{`RANDOM}};
  FifoCell_758 = _RAND_760[8:0];
  _RAND_761 = {1{`RANDOM}};
  FifoCell_759 = _RAND_761[8:0];
  _RAND_762 = {1{`RANDOM}};
  FifoCell_760 = _RAND_762[8:0];
  _RAND_763 = {1{`RANDOM}};
  FifoCell_761 = _RAND_763[8:0];
  _RAND_764 = {1{`RANDOM}};
  FifoCell_762 = _RAND_764[8:0];
  _RAND_765 = {1{`RANDOM}};
  FifoCell_763 = _RAND_765[8:0];
  _RAND_766 = {1{`RANDOM}};
  FifoCell_764 = _RAND_766[8:0];
  _RAND_767 = {1{`RANDOM}};
  FifoCell_765 = _RAND_767[8:0];
  _RAND_768 = {1{`RANDOM}};
  FifoCell_766 = _RAND_768[8:0];
  _RAND_769 = {1{`RANDOM}};
  FifoCell_767 = _RAND_769[8:0];
  _RAND_770 = {1{`RANDOM}};
  FifoCell_768 = _RAND_770[8:0];
  _RAND_771 = {1{`RANDOM}};
  FifoCell_769 = _RAND_771[8:0];
  _RAND_772 = {1{`RANDOM}};
  FifoCell_770 = _RAND_772[8:0];
  _RAND_773 = {1{`RANDOM}};
  FifoCell_771 = _RAND_773[8:0];
  _RAND_774 = {1{`RANDOM}};
  FifoCell_772 = _RAND_774[8:0];
  _RAND_775 = {1{`RANDOM}};
  FifoCell_773 = _RAND_775[8:0];
  _RAND_776 = {1{`RANDOM}};
  FifoCell_774 = _RAND_776[8:0];
  _RAND_777 = {1{`RANDOM}};
  FifoCell_775 = _RAND_777[8:0];
  _RAND_778 = {1{`RANDOM}};
  FifoCell_776 = _RAND_778[8:0];
  _RAND_779 = {1{`RANDOM}};
  FifoCell_777 = _RAND_779[8:0];
  _RAND_780 = {1{`RANDOM}};
  FifoCell_778 = _RAND_780[8:0];
  _RAND_781 = {1{`RANDOM}};
  FifoCell_779 = _RAND_781[8:0];
  _RAND_782 = {1{`RANDOM}};
  FifoCell_780 = _RAND_782[8:0];
  _RAND_783 = {1{`RANDOM}};
  FifoCell_781 = _RAND_783[8:0];
  _RAND_784 = {1{`RANDOM}};
  FifoCell_782 = _RAND_784[8:0];
  _RAND_785 = {1{`RANDOM}};
  FifoCell_783 = _RAND_785[8:0];
  _RAND_786 = {1{`RANDOM}};
  FifoCell_784 = _RAND_786[8:0];
  _RAND_787 = {1{`RANDOM}};
  FifoCell_785 = _RAND_787[8:0];
  _RAND_788 = {1{`RANDOM}};
  FifoCell_786 = _RAND_788[8:0];
  _RAND_789 = {1{`RANDOM}};
  FifoCell_787 = _RAND_789[8:0];
  _RAND_790 = {1{`RANDOM}};
  FifoCell_788 = _RAND_790[8:0];
  _RAND_791 = {1{`RANDOM}};
  FifoCell_789 = _RAND_791[8:0];
  _RAND_792 = {1{`RANDOM}};
  FifoCell_790 = _RAND_792[8:0];
  _RAND_793 = {1{`RANDOM}};
  FifoCell_791 = _RAND_793[8:0];
  _RAND_794 = {1{`RANDOM}};
  FifoCell_792 = _RAND_794[8:0];
  _RAND_795 = {1{`RANDOM}};
  FifoCell_793 = _RAND_795[8:0];
  _RAND_796 = {1{`RANDOM}};
  FifoCell_794 = _RAND_796[8:0];
  _RAND_797 = {1{`RANDOM}};
  FifoCell_795 = _RAND_797[8:0];
  _RAND_798 = {1{`RANDOM}};
  FifoCell_796 = _RAND_798[8:0];
  _RAND_799 = {1{`RANDOM}};
  FifoCell_797 = _RAND_799[8:0];
  _RAND_800 = {1{`RANDOM}};
  FifoCell_798 = _RAND_800[8:0];
  _RAND_801 = {1{`RANDOM}};
  FifoCell_799 = _RAND_801[8:0];
  _RAND_802 = {1{`RANDOM}};
  FifoCell_800 = _RAND_802[8:0];
  _RAND_803 = {1{`RANDOM}};
  FifoCell_801 = _RAND_803[8:0];
  _RAND_804 = {1{`RANDOM}};
  FifoCell_802 = _RAND_804[8:0];
  _RAND_805 = {1{`RANDOM}};
  FifoCell_803 = _RAND_805[8:0];
  _RAND_806 = {1{`RANDOM}};
  FifoCell_804 = _RAND_806[8:0];
  _RAND_807 = {1{`RANDOM}};
  FifoCell_805 = _RAND_807[8:0];
  _RAND_808 = {1{`RANDOM}};
  FifoCell_806 = _RAND_808[8:0];
  _RAND_809 = {1{`RANDOM}};
  FifoCell_807 = _RAND_809[8:0];
  _RAND_810 = {1{`RANDOM}};
  FifoCell_808 = _RAND_810[8:0];
  _RAND_811 = {1{`RANDOM}};
  FifoCell_809 = _RAND_811[8:0];
  _RAND_812 = {1{`RANDOM}};
  FifoCell_810 = _RAND_812[8:0];
  _RAND_813 = {1{`RANDOM}};
  FifoCell_811 = _RAND_813[8:0];
  _RAND_814 = {1{`RANDOM}};
  FifoCell_812 = _RAND_814[8:0];
  _RAND_815 = {1{`RANDOM}};
  FifoCell_813 = _RAND_815[8:0];
  _RAND_816 = {1{`RANDOM}};
  FifoCell_814 = _RAND_816[8:0];
  _RAND_817 = {1{`RANDOM}};
  FifoCell_815 = _RAND_817[8:0];
  _RAND_818 = {1{`RANDOM}};
  FifoCell_816 = _RAND_818[8:0];
  _RAND_819 = {1{`RANDOM}};
  FifoCell_817 = _RAND_819[8:0];
  _RAND_820 = {1{`RANDOM}};
  FifoCell_818 = _RAND_820[8:0];
  _RAND_821 = {1{`RANDOM}};
  FifoCell_819 = _RAND_821[8:0];
  _RAND_822 = {1{`RANDOM}};
  FifoCell_820 = _RAND_822[8:0];
  _RAND_823 = {1{`RANDOM}};
  FifoCell_821 = _RAND_823[8:0];
  _RAND_824 = {1{`RANDOM}};
  FifoCell_822 = _RAND_824[8:0];
  _RAND_825 = {1{`RANDOM}};
  FifoCell_823 = _RAND_825[8:0];
  _RAND_826 = {1{`RANDOM}};
  FifoCell_824 = _RAND_826[8:0];
  _RAND_827 = {1{`RANDOM}};
  FifoCell_825 = _RAND_827[8:0];
  _RAND_828 = {1{`RANDOM}};
  FifoCell_826 = _RAND_828[8:0];
  _RAND_829 = {1{`RANDOM}};
  FifoCell_827 = _RAND_829[8:0];
  _RAND_830 = {1{`RANDOM}};
  FifoCell_828 = _RAND_830[8:0];
  _RAND_831 = {1{`RANDOM}};
  FifoCell_829 = _RAND_831[8:0];
  _RAND_832 = {1{`RANDOM}};
  FifoCell_830 = _RAND_832[8:0];
  _RAND_833 = {1{`RANDOM}};
  FifoCell_831 = _RAND_833[8:0];
  _RAND_834 = {1{`RANDOM}};
  FifoCell_832 = _RAND_834[8:0];
  _RAND_835 = {1{`RANDOM}};
  FifoCell_833 = _RAND_835[8:0];
  _RAND_836 = {1{`RANDOM}};
  FifoCell_834 = _RAND_836[8:0];
  _RAND_837 = {1{`RANDOM}};
  FifoCell_835 = _RAND_837[8:0];
  _RAND_838 = {1{`RANDOM}};
  FifoCell_836 = _RAND_838[8:0];
  _RAND_839 = {1{`RANDOM}};
  FifoCell_837 = _RAND_839[8:0];
  _RAND_840 = {1{`RANDOM}};
  FifoCell_838 = _RAND_840[8:0];
  _RAND_841 = {1{`RANDOM}};
  FifoCell_839 = _RAND_841[8:0];
  _RAND_842 = {1{`RANDOM}};
  FifoCell_840 = _RAND_842[8:0];
  _RAND_843 = {1{`RANDOM}};
  FifoCell_841 = _RAND_843[8:0];
  _RAND_844 = {1{`RANDOM}};
  FifoCell_842 = _RAND_844[8:0];
  _RAND_845 = {1{`RANDOM}};
  FifoCell_843 = _RAND_845[8:0];
  _RAND_846 = {1{`RANDOM}};
  FifoCell_844 = _RAND_846[8:0];
  _RAND_847 = {1{`RANDOM}};
  FifoCell_845 = _RAND_847[8:0];
  _RAND_848 = {1{`RANDOM}};
  FifoCell_846 = _RAND_848[8:0];
  _RAND_849 = {1{`RANDOM}};
  FifoCell_847 = _RAND_849[8:0];
  _RAND_850 = {1{`RANDOM}};
  FifoCell_848 = _RAND_850[8:0];
  _RAND_851 = {1{`RANDOM}};
  FifoCell_849 = _RAND_851[8:0];
  _RAND_852 = {1{`RANDOM}};
  FifoCell_850 = _RAND_852[8:0];
  _RAND_853 = {1{`RANDOM}};
  FifoCell_851 = _RAND_853[8:0];
  _RAND_854 = {1{`RANDOM}};
  FifoCell_852 = _RAND_854[8:0];
  _RAND_855 = {1{`RANDOM}};
  FifoCell_853 = _RAND_855[8:0];
  _RAND_856 = {1{`RANDOM}};
  FifoCell_854 = _RAND_856[8:0];
  _RAND_857 = {1{`RANDOM}};
  FifoCell_855 = _RAND_857[8:0];
  _RAND_858 = {1{`RANDOM}};
  FifoCell_856 = _RAND_858[8:0];
  _RAND_859 = {1{`RANDOM}};
  FifoCell_857 = _RAND_859[8:0];
  _RAND_860 = {1{`RANDOM}};
  FifoCell_858 = _RAND_860[8:0];
  _RAND_861 = {1{`RANDOM}};
  FifoCell_859 = _RAND_861[8:0];
  _RAND_862 = {1{`RANDOM}};
  FifoCell_860 = _RAND_862[8:0];
  _RAND_863 = {1{`RANDOM}};
  FifoCell_861 = _RAND_863[8:0];
  _RAND_864 = {1{`RANDOM}};
  FifoCell_862 = _RAND_864[8:0];
  _RAND_865 = {1{`RANDOM}};
  FifoCell_863 = _RAND_865[8:0];
  _RAND_866 = {1{`RANDOM}};
  FifoCell_864 = _RAND_866[8:0];
  _RAND_867 = {1{`RANDOM}};
  FifoCell_865 = _RAND_867[8:0];
  _RAND_868 = {1{`RANDOM}};
  FifoCell_866 = _RAND_868[8:0];
  _RAND_869 = {1{`RANDOM}};
  FifoCell_867 = _RAND_869[8:0];
  _RAND_870 = {1{`RANDOM}};
  FifoCell_868 = _RAND_870[8:0];
  _RAND_871 = {1{`RANDOM}};
  FifoCell_869 = _RAND_871[8:0];
  _RAND_872 = {1{`RANDOM}};
  FifoCell_870 = _RAND_872[8:0];
  _RAND_873 = {1{`RANDOM}};
  FifoCell_871 = _RAND_873[8:0];
  _RAND_874 = {1{`RANDOM}};
  FifoCell_872 = _RAND_874[8:0];
  _RAND_875 = {1{`RANDOM}};
  FifoCell_873 = _RAND_875[8:0];
  _RAND_876 = {1{`RANDOM}};
  FifoCell_874 = _RAND_876[8:0];
  _RAND_877 = {1{`RANDOM}};
  FifoCell_875 = _RAND_877[8:0];
  _RAND_878 = {1{`RANDOM}};
  FifoCell_876 = _RAND_878[8:0];
  _RAND_879 = {1{`RANDOM}};
  FifoCell_877 = _RAND_879[8:0];
  _RAND_880 = {1{`RANDOM}};
  FifoCell_878 = _RAND_880[8:0];
  _RAND_881 = {1{`RANDOM}};
  FifoCell_879 = _RAND_881[8:0];
  _RAND_882 = {1{`RANDOM}};
  FifoCell_880 = _RAND_882[8:0];
  _RAND_883 = {1{`RANDOM}};
  FifoCell_881 = _RAND_883[8:0];
  _RAND_884 = {1{`RANDOM}};
  FifoCell_882 = _RAND_884[8:0];
  _RAND_885 = {1{`RANDOM}};
  FifoCell_883 = _RAND_885[8:0];
  _RAND_886 = {1{`RANDOM}};
  FifoCell_884 = _RAND_886[8:0];
  _RAND_887 = {1{`RANDOM}};
  FifoCell_885 = _RAND_887[8:0];
  _RAND_888 = {1{`RANDOM}};
  FifoCell_886 = _RAND_888[8:0];
  _RAND_889 = {1{`RANDOM}};
  FifoCell_887 = _RAND_889[8:0];
  _RAND_890 = {1{`RANDOM}};
  FifoCell_888 = _RAND_890[8:0];
  _RAND_891 = {1{`RANDOM}};
  FifoCell_889 = _RAND_891[8:0];
  _RAND_892 = {1{`RANDOM}};
  FifoCell_890 = _RAND_892[8:0];
  _RAND_893 = {1{`RANDOM}};
  FifoCell_891 = _RAND_893[8:0];
  _RAND_894 = {1{`RANDOM}};
  FifoCell_892 = _RAND_894[8:0];
  _RAND_895 = {1{`RANDOM}};
  FifoCell_893 = _RAND_895[8:0];
  _RAND_896 = {1{`RANDOM}};
  FifoCell_894 = _RAND_896[8:0];
  _RAND_897 = {1{`RANDOM}};
  FifoCell_895 = _RAND_897[8:0];
  _RAND_898 = {1{`RANDOM}};
  FifoCell_896 = _RAND_898[8:0];
  _RAND_899 = {1{`RANDOM}};
  FifoCell_897 = _RAND_899[8:0];
  _RAND_900 = {1{`RANDOM}};
  FifoCell_898 = _RAND_900[8:0];
  _RAND_901 = {1{`RANDOM}};
  FifoCell_899 = _RAND_901[8:0];
  _RAND_902 = {1{`RANDOM}};
  FifoCell_900 = _RAND_902[8:0];
  _RAND_903 = {1{`RANDOM}};
  FifoCell_901 = _RAND_903[8:0];
  _RAND_904 = {1{`RANDOM}};
  FifoCell_902 = _RAND_904[8:0];
  _RAND_905 = {1{`RANDOM}};
  FifoCell_903 = _RAND_905[8:0];
  _RAND_906 = {1{`RANDOM}};
  FifoCell_904 = _RAND_906[8:0];
  _RAND_907 = {1{`RANDOM}};
  FifoCell_905 = _RAND_907[8:0];
  _RAND_908 = {1{`RANDOM}};
  FifoCell_906 = _RAND_908[8:0];
  _RAND_909 = {1{`RANDOM}};
  FifoCell_907 = _RAND_909[8:0];
  _RAND_910 = {1{`RANDOM}};
  FifoCell_908 = _RAND_910[8:0];
  _RAND_911 = {1{`RANDOM}};
  FifoCell_909 = _RAND_911[8:0];
  _RAND_912 = {1{`RANDOM}};
  FifoCell_910 = _RAND_912[8:0];
  _RAND_913 = {1{`RANDOM}};
  FifoCell_911 = _RAND_913[8:0];
  _RAND_914 = {1{`RANDOM}};
  FifoCell_912 = _RAND_914[8:0];
  _RAND_915 = {1{`RANDOM}};
  FifoCell_913 = _RAND_915[8:0];
  _RAND_916 = {1{`RANDOM}};
  FifoCell_914 = _RAND_916[8:0];
  _RAND_917 = {1{`RANDOM}};
  FifoCell_915 = _RAND_917[8:0];
  _RAND_918 = {1{`RANDOM}};
  FifoCell_916 = _RAND_918[8:0];
  _RAND_919 = {1{`RANDOM}};
  FifoCell_917 = _RAND_919[8:0];
  _RAND_920 = {1{`RANDOM}};
  FifoCell_918 = _RAND_920[8:0];
  _RAND_921 = {1{`RANDOM}};
  FifoCell_919 = _RAND_921[8:0];
  _RAND_922 = {1{`RANDOM}};
  FifoCell_920 = _RAND_922[8:0];
  _RAND_923 = {1{`RANDOM}};
  FifoCell_921 = _RAND_923[8:0];
  _RAND_924 = {1{`RANDOM}};
  FifoCell_922 = _RAND_924[8:0];
  _RAND_925 = {1{`RANDOM}};
  FifoCell_923 = _RAND_925[8:0];
  _RAND_926 = {1{`RANDOM}};
  FifoCell_924 = _RAND_926[8:0];
  _RAND_927 = {1{`RANDOM}};
  FifoCell_925 = _RAND_927[8:0];
  _RAND_928 = {1{`RANDOM}};
  FifoCell_926 = _RAND_928[8:0];
  _RAND_929 = {1{`RANDOM}};
  FifoCell_927 = _RAND_929[8:0];
  _RAND_930 = {1{`RANDOM}};
  FifoCell_928 = _RAND_930[8:0];
  _RAND_931 = {1{`RANDOM}};
  FifoCell_929 = _RAND_931[8:0];
  _RAND_932 = {1{`RANDOM}};
  FifoCell_930 = _RAND_932[8:0];
  _RAND_933 = {1{`RANDOM}};
  FifoCell_931 = _RAND_933[8:0];
  _RAND_934 = {1{`RANDOM}};
  FifoCell_932 = _RAND_934[8:0];
  _RAND_935 = {1{`RANDOM}};
  FifoCell_933 = _RAND_935[8:0];
  _RAND_936 = {1{`RANDOM}};
  FifoCell_934 = _RAND_936[8:0];
  _RAND_937 = {1{`RANDOM}};
  FifoCell_935 = _RAND_937[8:0];
  _RAND_938 = {1{`RANDOM}};
  FifoCell_936 = _RAND_938[8:0];
  _RAND_939 = {1{`RANDOM}};
  FifoCell_937 = _RAND_939[8:0];
  _RAND_940 = {1{`RANDOM}};
  FifoCell_938 = _RAND_940[8:0];
  _RAND_941 = {1{`RANDOM}};
  FifoCell_939 = _RAND_941[8:0];
  _RAND_942 = {1{`RANDOM}};
  FifoCell_940 = _RAND_942[8:0];
  _RAND_943 = {1{`RANDOM}};
  FifoCell_941 = _RAND_943[8:0];
  _RAND_944 = {1{`RANDOM}};
  FifoCell_942 = _RAND_944[8:0];
  _RAND_945 = {1{`RANDOM}};
  FifoCell_943 = _RAND_945[8:0];
  _RAND_946 = {1{`RANDOM}};
  FifoCell_944 = _RAND_946[8:0];
  _RAND_947 = {1{`RANDOM}};
  FifoCell_945 = _RAND_947[8:0];
  _RAND_948 = {1{`RANDOM}};
  FifoCell_946 = _RAND_948[8:0];
  _RAND_949 = {1{`RANDOM}};
  FifoCell_947 = _RAND_949[8:0];
  _RAND_950 = {1{`RANDOM}};
  FifoCell_948 = _RAND_950[8:0];
  _RAND_951 = {1{`RANDOM}};
  FifoCell_949 = _RAND_951[8:0];
  _RAND_952 = {1{`RANDOM}};
  FifoCell_950 = _RAND_952[8:0];
  _RAND_953 = {1{`RANDOM}};
  FifoCell_951 = _RAND_953[8:0];
  _RAND_954 = {1{`RANDOM}};
  FifoCell_952 = _RAND_954[8:0];
  _RAND_955 = {1{`RANDOM}};
  FifoCell_953 = _RAND_955[8:0];
  _RAND_956 = {1{`RANDOM}};
  FifoCell_954 = _RAND_956[8:0];
  _RAND_957 = {1{`RANDOM}};
  FifoCell_955 = _RAND_957[8:0];
  _RAND_958 = {1{`RANDOM}};
  FifoCell_956 = _RAND_958[8:0];
  _RAND_959 = {1{`RANDOM}};
  FifoCell_957 = _RAND_959[8:0];
  _RAND_960 = {1{`RANDOM}};
  FifoCell_958 = _RAND_960[8:0];
  _RAND_961 = {1{`RANDOM}};
  FifoCell_959 = _RAND_961[8:0];
  _RAND_962 = {1{`RANDOM}};
  FifoCell_960 = _RAND_962[8:0];
  _RAND_963 = {1{`RANDOM}};
  FifoCell_961 = _RAND_963[8:0];
  _RAND_964 = {1{`RANDOM}};
  FifoCell_962 = _RAND_964[8:0];
  _RAND_965 = {1{`RANDOM}};
  FifoCell_963 = _RAND_965[8:0];
  _RAND_966 = {1{`RANDOM}};
  FifoCell_964 = _RAND_966[8:0];
  _RAND_967 = {1{`RANDOM}};
  FifoCell_965 = _RAND_967[8:0];
  _RAND_968 = {1{`RANDOM}};
  FifoCell_966 = _RAND_968[8:0];
  _RAND_969 = {1{`RANDOM}};
  FifoCell_967 = _RAND_969[8:0];
  _RAND_970 = {1{`RANDOM}};
  FifoCell_968 = _RAND_970[8:0];
  _RAND_971 = {1{`RANDOM}};
  FifoCell_969 = _RAND_971[8:0];
  _RAND_972 = {1{`RANDOM}};
  FifoCell_970 = _RAND_972[8:0];
  _RAND_973 = {1{`RANDOM}};
  FifoCell_971 = _RAND_973[8:0];
  _RAND_974 = {1{`RANDOM}};
  FifoCell_972 = _RAND_974[8:0];
  _RAND_975 = {1{`RANDOM}};
  FifoCell_973 = _RAND_975[8:0];
  _RAND_976 = {1{`RANDOM}};
  FifoCell_974 = _RAND_976[8:0];
  _RAND_977 = {1{`RANDOM}};
  FifoCell_975 = _RAND_977[8:0];
  _RAND_978 = {1{`RANDOM}};
  FifoCell_976 = _RAND_978[8:0];
  _RAND_979 = {1{`RANDOM}};
  FifoCell_977 = _RAND_979[8:0];
  _RAND_980 = {1{`RANDOM}};
  FifoCell_978 = _RAND_980[8:0];
  _RAND_981 = {1{`RANDOM}};
  FifoCell_979 = _RAND_981[8:0];
  _RAND_982 = {1{`RANDOM}};
  FifoCell_980 = _RAND_982[8:0];
  _RAND_983 = {1{`RANDOM}};
  FifoCell_981 = _RAND_983[8:0];
  _RAND_984 = {1{`RANDOM}};
  FifoCell_982 = _RAND_984[8:0];
  _RAND_985 = {1{`RANDOM}};
  FifoCell_983 = _RAND_985[8:0];
  _RAND_986 = {1{`RANDOM}};
  FifoCell_984 = _RAND_986[8:0];
  _RAND_987 = {1{`RANDOM}};
  FifoCell_985 = _RAND_987[8:0];
  _RAND_988 = {1{`RANDOM}};
  FifoCell_986 = _RAND_988[8:0];
  _RAND_989 = {1{`RANDOM}};
  FifoCell_987 = _RAND_989[8:0];
  _RAND_990 = {1{`RANDOM}};
  FifoCell_988 = _RAND_990[8:0];
  _RAND_991 = {1{`RANDOM}};
  FifoCell_989 = _RAND_991[8:0];
  _RAND_992 = {1{`RANDOM}};
  FifoCell_990 = _RAND_992[8:0];
  _RAND_993 = {1{`RANDOM}};
  FifoCell_991 = _RAND_993[8:0];
  _RAND_994 = {1{`RANDOM}};
  FifoCell_992 = _RAND_994[8:0];
  _RAND_995 = {1{`RANDOM}};
  FifoCell_993 = _RAND_995[8:0];
  _RAND_996 = {1{`RANDOM}};
  FifoCell_994 = _RAND_996[8:0];
  _RAND_997 = {1{`RANDOM}};
  FifoCell_995 = _RAND_997[8:0];
  _RAND_998 = {1{`RANDOM}};
  FifoCell_996 = _RAND_998[8:0];
  _RAND_999 = {1{`RANDOM}};
  FifoCell_997 = _RAND_999[8:0];
  _RAND_1000 = {1{`RANDOM}};
  FifoCell_998 = _RAND_1000[8:0];
  _RAND_1001 = {1{`RANDOM}};
  FifoCell_999 = _RAND_1001[8:0];
  _RAND_1002 = {1{`RANDOM}};
  FifoCell_1000 = _RAND_1002[8:0];
  _RAND_1003 = {1{`RANDOM}};
  FifoCell_1001 = _RAND_1003[8:0];
  _RAND_1004 = {1{`RANDOM}};
  FifoCell_1002 = _RAND_1004[8:0];
  _RAND_1005 = {1{`RANDOM}};
  FifoCell_1003 = _RAND_1005[8:0];
  _RAND_1006 = {1{`RANDOM}};
  FifoCell_1004 = _RAND_1006[8:0];
  _RAND_1007 = {1{`RANDOM}};
  FifoCell_1005 = _RAND_1007[8:0];
  _RAND_1008 = {1{`RANDOM}};
  FifoCell_1006 = _RAND_1008[8:0];
  _RAND_1009 = {1{`RANDOM}};
  FifoCell_1007 = _RAND_1009[8:0];
  _RAND_1010 = {1{`RANDOM}};
  FifoCell_1008 = _RAND_1010[8:0];
  _RAND_1011 = {1{`RANDOM}};
  FifoCell_1009 = _RAND_1011[8:0];
  _RAND_1012 = {1{`RANDOM}};
  FifoCell_1010 = _RAND_1012[8:0];
  _RAND_1013 = {1{`RANDOM}};
  FifoCell_1011 = _RAND_1013[8:0];
  _RAND_1014 = {1{`RANDOM}};
  FifoCell_1012 = _RAND_1014[8:0];
  _RAND_1015 = {1{`RANDOM}};
  FifoCell_1013 = _RAND_1015[8:0];
  _RAND_1016 = {1{`RANDOM}};
  FifoCell_1014 = _RAND_1016[8:0];
  _RAND_1017 = {1{`RANDOM}};
  FifoCell_1015 = _RAND_1017[8:0];
  _RAND_1018 = {1{`RANDOM}};
  FifoCell_1016 = _RAND_1018[8:0];
  _RAND_1019 = {1{`RANDOM}};
  FifoCell_1017 = _RAND_1019[8:0];
  _RAND_1020 = {1{`RANDOM}};
  FifoCell_1018 = _RAND_1020[8:0];
  _RAND_1021 = {1{`RANDOM}};
  FifoCell_1019 = _RAND_1021[8:0];
  _RAND_1022 = {1{`RANDOM}};
  FifoCell_1020 = _RAND_1022[8:0];
  _RAND_1023 = {1{`RANDOM}};
  FifoCell_1021 = _RAND_1023[8:0];
  _RAND_1024 = {1{`RANDOM}};
  FifoCell_1022 = _RAND_1024[8:0];
  _RAND_1025 = {1{`RANDOM}};
  FifoCell_1023 = _RAND_1025[8:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module AxisCrcChecker(
  input        clock,
  input        reset,
  output       io_AxisSlv_ready, // @[src/main/scala/axis_crc_ckecker_pkg/AxisCrcChecker.scala 23:14]
  input        io_AxisSlv_valid, // @[src/main/scala/axis_crc_ckecker_pkg/AxisCrcChecker.scala 23:14]
  input        io_AxisSlv_bits_Tlast, // @[src/main/scala/axis_crc_ckecker_pkg/AxisCrcChecker.scala 23:14]
  input  [7:0] io_AxisSlv_bits_Tdata, // @[src/main/scala/axis_crc_ckecker_pkg/AxisCrcChecker.scala 23:14]
  input        io_AxisMst_ready, // @[src/main/scala/axis_crc_ckecker_pkg/AxisCrcChecker.scala 23:14]
  output       io_AxisMst_valid, // @[src/main/scala/axis_crc_ckecker_pkg/AxisCrcChecker.scala 23:14]
  output       io_AxisMst_bits_Tlast, // @[src/main/scala/axis_crc_ckecker_pkg/AxisCrcChecker.scala 23:14]
  output [7:0] io_AxisMst_bits_Tdata // @[src/main/scala/axis_crc_ckecker_pkg/AxisCrcChecker.scala 23:14]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  wire [7:0] u_calc_crc_CRC_I; // @[src/main/scala/axis_crc_ckecker_pkg/AxisCrcChecker.scala 85:26]
  wire [7:0] u_calc_crc_DATA_I; // @[src/main/scala/axis_crc_ckecker_pkg/AxisCrcChecker.scala 85:26]
  wire [7:0] u_calc_crc_CRC_O; // @[src/main/scala/axis_crc_ckecker_pkg/AxisCrcChecker.scala 85:26]
  wire  u_sync_fifo_clock; // @[src/main/scala/axis_crc_ckecker_pkg/AxisCrcChecker.scala 93:27]
  wire  u_sync_fifo_reset; // @[src/main/scala/axis_crc_ckecker_pkg/AxisCrcChecker.scala 93:27]
  wire  u_sync_fifo_io_Writer_WriteEn; // @[src/main/scala/axis_crc_ckecker_pkg/AxisCrcChecker.scala 93:27]
  wire [8:0] u_sync_fifo_io_Writer_WriteData; // @[src/main/scala/axis_crc_ckecker_pkg/AxisCrcChecker.scala 93:27]
  wire  u_sync_fifo_io_Writer_Full; // @[src/main/scala/axis_crc_ckecker_pkg/AxisCrcChecker.scala 93:27]
  wire  u_sync_fifo_io_Reader_ReadEn; // @[src/main/scala/axis_crc_ckecker_pkg/AxisCrcChecker.scala 93:27]
  wire [8:0] u_sync_fifo_io_Reader_ReadData; // @[src/main/scala/axis_crc_ckecker_pkg/AxisCrcChecker.scala 93:27]
  wire  u_sync_fifo_io_Reader_Empty; // @[src/main/scala/axis_crc_ckecker_pkg/AxisCrcChecker.scala 93:27]
  reg [7:0] CrcInReg; // @[src/main/scala/axis_crc_ckecker_pkg/AxisCrcChecker.scala 30:32]
  reg  FifoRstReg; // @[src/main/scala/axis_crc_ckecker_pkg/AxisCrcChecker.scala 32:32]
  reg [1:0] CheckerStReg; // @[src/main/scala/axis_crc_ckecker_pkg/AxisCrcChecker.scala 38:29]
  wire  _PacketReceived_T = io_AxisSlv_valid & io_AxisSlv_ready; // @[src/main/scala/axis_crc_ckecker_pkg/AxisCrcChecker.scala 40:38]
  wire  PacketReceived = io_AxisSlv_valid & io_AxisSlv_ready & io_AxisSlv_bits_Tlast; // @[src/main/scala/axis_crc_ckecker_pkg/AxisCrcChecker.scala 40:57]
  wire  RacketSended = io_AxisMst_valid & io_AxisMst_ready & io_AxisMst_bits_Tlast; // @[src/main/scala/axis_crc_ckecker_pkg/AxisCrcChecker.scala 42:55]
  wire [1:0] _GEN_2 = RacketSended ? 2'h0 : CheckerStReg; // @[src/main/scala/axis_crc_ckecker_pkg/AxisCrcChecker.scala 62:35 63:22 38:29]
  wire [1:0] _GEN_3 = 2'h3 == CheckerStReg ? _GEN_2 : CheckerStReg; // @[src/main/scala/axis_crc_ckecker_pkg/AxisCrcChecker.scala 44:25 38:29]
  reg  AxisSlvTready; // @[src/main/scala/axis_crc_ckecker_pkg/AxisCrcChecker.scala 68:30]
  wire  _GEN_7 = CheckerStReg == 2'h0 | AxisSlvTready; // @[src/main/scala/axis_crc_ckecker_pkg/AxisCrcChecker.scala 72:43 73:19 68:30]
  wire [7:0] CrcOut = u_calc_crc_CRC_O; // @[src/main/scala/axis_crc_ckecker_pkg/AxisCrcChecker.scala 31:29 89:25]
  wire  _u_sync_fifo_io_Reader_ReadEn_T = CheckerStReg == 2'h3; // @[src/main/scala/axis_crc_ckecker_pkg/AxisCrcChecker.scala 100:49]
  calc_crc u_calc_crc ( // @[src/main/scala/axis_crc_ckecker_pkg/AxisCrcChecker.scala 85:26]
    .CRC_I(u_calc_crc_CRC_I),
    .DATA_I(u_calc_crc_DATA_I),
    .CRC_O(u_calc_crc_CRC_O)
  );
  SyncFifo u_sync_fifo ( // @[src/main/scala/axis_crc_ckecker_pkg/AxisCrcChecker.scala 93:27]
    .clock(u_sync_fifo_clock),
    .reset(u_sync_fifo_reset),
    .io_Writer_WriteEn(u_sync_fifo_io_Writer_WriteEn),
    .io_Writer_WriteData(u_sync_fifo_io_Writer_WriteData),
    .io_Writer_Full(u_sync_fifo_io_Writer_Full),
    .io_Reader_ReadEn(u_sync_fifo_io_Reader_ReadEn),
    .io_Reader_ReadData(u_sync_fifo_io_Reader_ReadData),
    .io_Reader_Empty(u_sync_fifo_io_Reader_Empty)
  );
  assign io_AxisSlv_ready = AxisSlvTready; // @[src/main/scala/axis_crc_ckecker_pkg/AxisCrcChecker.scala 76:20]
  assign io_AxisMst_valid = _u_sync_fifo_io_Reader_ReadEn_T & ~u_sync_fifo_io_Reader_Empty; // @[src/main/scala/axis_crc_ckecker_pkg/AxisCrcChecker.scala 102:49]
  assign io_AxisMst_bits_Tlast = u_sync_fifo_io_Reader_ReadData[8]; // @[src/main/scala/axis_crc_ckecker_pkg/AxisCrcChecker.scala 105:58]
  assign io_AxisMst_bits_Tdata = u_sync_fifo_io_Reader_ReadData[7:0]; // @[src/main/scala/axis_crc_ckecker_pkg/AxisCrcChecker.scala 104:58]
  assign u_calc_crc_CRC_I = CrcInReg; // @[src/main/scala/axis_crc_ckecker_pkg/AxisCrcChecker.scala 87:25]
  assign u_calc_crc_DATA_I = io_AxisSlv_bits_Tdata; // @[src/main/scala/axis_crc_ckecker_pkg/AxisCrcChecker.scala 88:25]
  assign u_sync_fifo_clock = clock;
  assign u_sync_fifo_reset = FifoRstReg; // @[src/main/scala/axis_crc_ckecker_pkg/AxisCrcChecker.scala 95:36]
  assign u_sync_fifo_io_Writer_WriteEn = io_AxisSlv_valid & io_AxisSlv_ready; // @[src/main/scala/axis_crc_ckecker_pkg/AxisCrcChecker.scala 98:53]
  assign u_sync_fifo_io_Writer_WriteData = {io_AxisSlv_bits_Tlast,io_AxisSlv_bits_Tdata}; // @[src/main/scala/axis_crc_ckecker_pkg/AxisCrcChecker.scala 97:60]
  assign u_sync_fifo_io_Reader_ReadEn = CheckerStReg == 2'h3 & io_AxisMst_ready; // @[src/main/scala/axis_crc_ckecker_pkg/AxisCrcChecker.scala 100:61]
  always @(posedge clock) begin
    if (reset) begin // @[src/main/scala/axis_crc_ckecker_pkg/AxisCrcChecker.scala 30:32]
      CrcInReg <= 8'hff; // @[src/main/scala/axis_crc_ckecker_pkg/AxisCrcChecker.scala 30:32]
    end else if (_PacketReceived_T) begin // @[src/main/scala/axis_crc_ckecker_pkg/AxisCrcChecker.scala 78:46]
      CrcInReg <= CrcOut; // @[src/main/scala/axis_crc_ckecker_pkg/AxisCrcChecker.scala 79:14]
    end else if (CheckerStReg == 2'h1) begin // @[src/main/scala/axis_crc_ckecker_pkg/AxisCrcChecker.scala 81:41]
      CrcInReg <= 8'hff; // @[src/main/scala/axis_crc_ckecker_pkg/AxisCrcChecker.scala 82:14]
    end
    FifoRstReg <= reset | CheckerStReg == 2'h2; // @[src/main/scala/axis_crc_ckecker_pkg/AxisCrcChecker.scala 32:{32,32} 91:14]
    if (reset) begin // @[src/main/scala/axis_crc_ckecker_pkg/AxisCrcChecker.scala 38:29]
      CheckerStReg <= 2'h0; // @[src/main/scala/axis_crc_ckecker_pkg/AxisCrcChecker.scala 38:29]
    end else if (2'h0 == CheckerStReg) begin // @[src/main/scala/axis_crc_ckecker_pkg/AxisCrcChecker.scala 44:25]
      if (PacketReceived) begin // @[src/main/scala/axis_crc_ckecker_pkg/AxisCrcChecker.scala 46:37]
        CheckerStReg <= 2'h1; // @[src/main/scala/axis_crc_ckecker_pkg/AxisCrcChecker.scala 47:22]
      end
    end else if (2'h1 == CheckerStReg) begin // @[src/main/scala/axis_crc_ckecker_pkg/AxisCrcChecker.scala 44:25]
      if (CrcInReg == 8'h0) begin // @[src/main/scala/axis_crc_ckecker_pkg/AxisCrcChecker.scala 51:31]
        CheckerStReg <= 2'h3; // @[src/main/scala/axis_crc_ckecker_pkg/AxisCrcChecker.scala 52:22]
      end else begin
        CheckerStReg <= 2'h2; // @[src/main/scala/axis_crc_ckecker_pkg/AxisCrcChecker.scala 55:22]
      end
    end else if (2'h2 == CheckerStReg) begin // @[src/main/scala/axis_crc_ckecker_pkg/AxisCrcChecker.scala 44:25]
      CheckerStReg <= 2'h0; // @[src/main/scala/axis_crc_ckecker_pkg/AxisCrcChecker.scala 59:20]
    end else begin
      CheckerStReg <= _GEN_3;
    end
    if (reset) begin // @[src/main/scala/axis_crc_ckecker_pkg/AxisCrcChecker.scala 68:30]
      AxisSlvTready <= 1'h0; // @[src/main/scala/axis_crc_ckecker_pkg/AxisCrcChecker.scala 68:30]
    end else if (PacketReceived) begin // @[src/main/scala/axis_crc_ckecker_pkg/AxisCrcChecker.scala 69:33]
      AxisSlvTready <= 1'h0; // @[src/main/scala/axis_crc_ckecker_pkg/AxisCrcChecker.scala 70:19]
    end else begin
      AxisSlvTready <= _GEN_7;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  CrcInReg = _RAND_0[7:0];
  _RAND_1 = {1{`RANDOM}};
  FifoRstReg = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  CheckerStReg = _RAND_2[1:0];
  _RAND_3 = {1{`RANDOM}};
  AxisSlvTready = _RAND_3[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
